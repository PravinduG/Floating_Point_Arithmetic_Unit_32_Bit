`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11/27/2025 09:45:09 PM
// Design Name: 
// Module Name: reciprocal_lut
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module reciprocal_lut(
			 input logic  [9:0]														lut_idx
			,output logic [31:0]													X0

    );
		
		always_comb begin
    case(lut_idx)
        10'd0 : X0 <= 32'h80000000;
        10'd1 : X0 <= 32'h7FE007FE;
        10'd2 : X0 <= 32'h7FC01FF0;
        10'd3 : X0 <= 32'h7FA047CA;
        10'd4 : X0 <= 32'h7F807F80;
        10'd5 : X0 <= 32'h7F60C707;
        10'd6 : X0 <= 32'h7F411E53;
        10'd7 : X0 <= 32'h7F218557;
        10'd8 : X0 <= 32'h7F01FC08;
        10'd9 : X0 <= 32'h7EE2825B;
        10'd10 : X0 <= 32'h7EC31843;
        10'd11 : X0 <= 32'h7EA3BDB6;
        10'd12 : X0 <= 32'h7E8472A8;
        10'd13 : X0 <= 32'h7E65370D;
        10'd14 : X0 <= 32'h7E460ADA;
        10'd15 : X0 <= 32'h7E26EE03;
        10'd16 : X0 <= 32'h7E07E07E;
        10'd17 : X0 <= 32'h7DE8E23E;
        10'd18 : X0 <= 32'h7DC9F339;
        10'd19 : X0 <= 32'h7DAB1364;
        10'd20 : X0 <= 32'h7D8C42B3;
        10'd21 : X0 <= 32'h7D6D811A;
        10'd22 : X0 <= 32'h7D4ECE90;
        10'd23 : X0 <= 32'h7D302B09;
        10'd24 : X0 <= 32'h7D119679;
        10'd25 : X0 <= 32'h7CF310D7;
        10'd26 : X0 <= 32'h7CD49A16;
        10'd27 : X0 <= 32'h7CB6322D;
        10'd28 : X0 <= 32'h7C97D911;
        10'd29 : X0 <= 32'h7C798EB5;
        10'd30 : X0 <= 32'h7C5B5311;
        10'd31 : X0 <= 32'h7C3D2619;
        10'd32 : X0 <= 32'h7C1F07C2;
        10'd33 : X0 <= 32'h7C00F802;
        10'd34 : X0 <= 32'h7BE2F6CE;
        10'd35 : X0 <= 32'h7BC5041C;
        10'd36 : X0 <= 32'h7BA71FE1;
        10'd37 : X0 <= 32'h7B894A13;
        10'd38 : X0 <= 32'h7B6B82A7;
        10'd39 : X0 <= 32'h7B4DC993;
        10'd40 : X0 <= 32'h7B301ECC;
        10'd41 : X0 <= 32'h7B128249;
        10'd42 : X0 <= 32'h7AF4F3FE;
        10'd43 : X0 <= 32'h7AD773E2;
        10'd44 : X0 <= 32'h7ABA01EB;
        10'd45 : X0 <= 32'h7A9C9E0E;
        10'd46 : X0 <= 32'h7A7F4841;
        10'd47 : X0 <= 32'h7A62007A;
        10'd48 : X0 <= 32'h7A44C6B0;
        10'd49 : X0 <= 32'h7A279AD7;
        10'd50 : X0 <= 32'h7A0A7CE7;
        10'd51 : X0 <= 32'h79ED6CD4;
        10'd52 : X0 <= 32'h79D06A96;
        10'd53 : X0 <= 32'h79B37623;
        10'd54 : X0 <= 32'h79968F70;
        10'd55 : X0 <= 32'h7979B673;
        10'd56 : X0 <= 32'h795CEB24;
        10'd57 : X0 <= 32'h79402D78;
        10'd58 : X0 <= 32'h79237D66;
        10'd59 : X0 <= 32'h7906DAE3;
        10'd60 : X0 <= 32'h78EA45E7;
        10'd61 : X0 <= 32'h78CDBE68;
        10'd62 : X0 <= 32'h78B1445C;
        10'd63 : X0 <= 32'h7894D7BA;
        10'd64 : X0 <= 32'h78787878;
        10'd65 : X0 <= 32'h785C268E;
        10'd66 : X0 <= 32'h783FE1F0;
        10'd67 : X0 <= 32'h7823AA97;
        10'd68 : X0 <= 32'h78078078;
        10'd69 : X0 <= 32'h77EB638B;
        10'd70 : X0 <= 32'h77CF53C6;
        10'd71 : X0 <= 32'h77B35120;
        10'd72 : X0 <= 32'h77975B90;
        10'd73 : X0 <= 32'h777B730C;
        10'd74 : X0 <= 32'h775F978C;
        10'd75 : X0 <= 32'h7743C907;
        10'd76 : X0 <= 32'h77280773;
        10'd77 : X0 <= 32'h770C52C7;
        10'd78 : X0 <= 32'h76F0AAFA;
        10'd79 : X0 <= 32'h76D51004;
        10'd80 : X0 <= 32'h76B981DB;
        10'd81 : X0 <= 32'h769E0077;
        10'd82 : X0 <= 32'h76828BCE;
        10'd83 : X0 <= 32'h766723D8;
        10'd84 : X0 <= 32'h764BC88C;
        10'd85 : X0 <= 32'h763079E2;
        10'd86 : X0 <= 32'h761537D0;
        10'd87 : X0 <= 32'h75FA024E;
        10'd88 : X0 <= 32'h75DED953;
        10'd89 : X0 <= 32'h75C3BCD6;
        10'd90 : X0 <= 32'h75A8ACD0;
        10'd91 : X0 <= 32'h758DA936;
        10'd92 : X0 <= 32'h7572B202;
        10'd93 : X0 <= 32'h7557C729;
        10'd94 : X0 <= 32'h753CE8A5;
        10'd95 : X0 <= 32'h7522166C;
        10'd96 : X0 <= 32'h75075075;
        10'd97 : X0 <= 32'h74EC96B9;
        10'd98 : X0 <= 32'h74D1E92F;
        10'd99 : X0 <= 32'h74B747CF;
        10'd100 : X0 <= 32'h749CB290;
        10'd101 : X0 <= 32'h7482296A;
        10'd102 : X0 <= 32'h7467AC55;
        10'd103 : X0 <= 32'h744D3B49;
        10'd104 : X0 <= 32'h7432D63E;
        10'd105 : X0 <= 32'h74187D2A;
        10'd106 : X0 <= 32'h73FE3007;
        10'd107 : X0 <= 32'h73E3EECC;
        10'd108 : X0 <= 32'h73C9B971;
        10'd109 : X0 <= 32'h73AF8FEE;
        10'd110 : X0 <= 32'h7395723B;
        10'd111 : X0 <= 32'h737B604F;
        10'd112 : X0 <= 32'h73615A24;
        10'd113 : X0 <= 32'h73475FB1;
        10'd114 : X0 <= 32'h732D70EE;
        10'd115 : X0 <= 32'h73138DD3;
        10'd116 : X0 <= 32'h72F9B658;
        10'd117 : X0 <= 32'h72DFEA76;
        10'd118 : X0 <= 32'h72C62A25;
        10'd119 : X0 <= 32'h72AC755D;
        10'd120 : X0 <= 32'h7292CC15;
        10'd121 : X0 <= 32'h72792E48;
        10'd122 : X0 <= 32'h725F9BEC;
        10'd123 : X0 <= 32'h724614FB;
        10'd124 : X0 <= 32'h722C996C;
        10'd125 : X0 <= 32'h72132938;
        10'd126 : X0 <= 32'h71F9C457;
        10'd127 : X0 <= 32'h71E06AC2;
        10'd128 : X0 <= 32'h71C71C72;
        10'd129 : X0 <= 32'h71ADD95E;
        10'd130 : X0 <= 32'h7194A17F;
        10'd131 : X0 <= 32'h717B74CF;
        10'd132 : X0 <= 32'h71625344;
        10'd133 : X0 <= 32'h71493CD9;
        10'd134 : X0 <= 32'h71303185;
        10'd135 : X0 <= 32'h71173142;
        10'd136 : X0 <= 32'h70FE3C07;
        10'd137 : X0 <= 32'h70E551CE;
        10'd138 : X0 <= 32'h70CC7290;
        10'd139 : X0 <= 32'h70B39E44;
        10'd140 : X0 <= 32'h709AD4E5;
        10'd141 : X0 <= 32'h7082166A;
        10'd142 : X0 <= 32'h706962CD;
        10'd143 : X0 <= 32'h7050BA06;
        10'd144 : X0 <= 32'h70381C0E;
        10'd145 : X0 <= 32'h701F88DE;
        10'd146 : X0 <= 32'h70070070;
        10'd147 : X0 <= 32'h6FEE82BC;
        10'd148 : X0 <= 32'h6FD60FBA;
        10'd149 : X0 <= 32'h6FBDA765;
        10'd150 : X0 <= 32'h6FA549B4;
        10'd151 : X0 <= 32'h6F8CF6A2;
        10'd152 : X0 <= 32'h6F74AE26;
        10'd153 : X0 <= 32'h6F5C703B;
        10'd154 : X0 <= 32'h6F443CD9;
        10'd155 : X0 <= 32'h6F2C13FA;
        10'd156 : X0 <= 32'h6F13F596;
        10'd157 : X0 <= 32'h6EFBE1A7;
        10'd158 : X0 <= 32'h6EE3D826;
        10'd159 : X0 <= 32'h6ECBD90C;
        10'd160 : X0 <= 32'h6EB3E453;
        10'd161 : X0 <= 32'h6E9BF9F3;
        10'd162 : X0 <= 32'h6E8419E7;
        10'd163 : X0 <= 32'h6E6C4427;
        10'd164 : X0 <= 32'h6E5478AC;
        10'd165 : X0 <= 32'h6E3CB771;
        10'd166 : X0 <= 32'h6E25006E;
        10'd167 : X0 <= 32'h6E0D539D;
        10'd168 : X0 <= 32'h6DF5B0F7;
        10'd169 : X0 <= 32'h6DDE1876;
        10'd170 : X0 <= 32'h6DC68A14;
        10'd171 : X0 <= 32'h6DAF05C9;
        10'd172 : X0 <= 32'h6D978B8F;
        10'd173 : X0 <= 32'h6D801B60;
        10'd174 : X0 <= 32'h6D68B535;
        10'd175 : X0 <= 32'h6D515909;
        10'd176 : X0 <= 32'h6D3A06D4;
        10'd177 : X0 <= 32'h6D22BE90;
        10'd178 : X0 <= 32'h6D0B8037;
        10'd179 : X0 <= 32'h6CF44BC2;
        10'd180 : X0 <= 32'h6CDD212B;
        10'd181 : X0 <= 32'h6CC6006D;
        10'd182 : X0 <= 32'h6CAEE980;
        10'd183 : X0 <= 32'h6C97DC5E;
        10'd184 : X0 <= 32'h6C80D902;
        10'd185 : X0 <= 32'h6C69DF64;
        10'd186 : X0 <= 32'h6C52EF7F;
        10'd187 : X0 <= 32'h6C3C094D;
        10'd188 : X0 <= 32'h6C252CC7;
        10'd189 : X0 <= 32'h6C0E59E8;
        10'd190 : X0 <= 32'h6BF790A9;
        10'd191 : X0 <= 32'h6BE0D104;
        10'd192 : X0 <= 32'h6BCA1AF3;
        10'd193 : X0 <= 32'h6BB36E6F;
        10'd194 : X0 <= 32'h6B9CCB74;
        10'd195 : X0 <= 32'h6B8631FB;
        10'd196 : X0 <= 32'h6B6FA1FE;
        10'd197 : X0 <= 32'h6B591B77;
        10'd198 : X0 <= 32'h6B429E60;
        10'd199 : X0 <= 32'h6B2C2AB4;
        10'd200 : X0 <= 32'h6B15C06B;
        10'd201 : X0 <= 32'h6AFF5F81;
        10'd202 : X0 <= 32'h6AE907EF;
        10'd203 : X0 <= 32'h6AD2B9B0;
        10'd204 : X0 <= 32'h6ABC74BE;
        10'd205 : X0 <= 32'h6AA63913;
        10'd206 : X0 <= 32'h6A9006A9;
        10'd207 : X0 <= 32'h6A79DD7A;
        10'd208 : X0 <= 32'h6A63BD82;
        10'd209 : X0 <= 32'h6A4DA6B9;
        10'd210 : X0 <= 32'h6A37991A;
        10'd211 : X0 <= 32'h6A2194A0;
        10'd212 : X0 <= 32'h6A0B9945;
        10'd213 : X0 <= 32'h69F5A703;
        10'd214 : X0 <= 32'h69DFBDD4;
        10'd215 : X0 <= 32'h69C9DDB4;
        10'd216 : X0 <= 32'h69B4069B;
        10'd217 : X0 <= 32'h699E3886;
        10'd218 : X0 <= 32'h6988736D;
        10'd219 : X0 <= 32'h6972B74C;
        10'd220 : X0 <= 32'h695D041E;
        10'd221 : X0 <= 32'h694759DB;
        10'd222 : X0 <= 32'h6931B880;
        10'd223 : X0 <= 32'h691C2007;
        10'd224 : X0 <= 32'h69069069;
        10'd225 : X0 <= 32'h68F109A2;
        10'd226 : X0 <= 32'h68DB8BAC;
        10'd227 : X0 <= 32'h68C61683;
        10'd228 : X0 <= 32'h68B0AA1F;
        10'd229 : X0 <= 32'h689B467D;
        10'd230 : X0 <= 32'h6885EB96;
        10'd231 : X0 <= 32'h68709965;
        10'd232 : X0 <= 32'h685B4FE6;
        10'd233 : X0 <= 32'h68460F12;
        10'd234 : X0 <= 32'h6830D6E5;
        10'd235 : X0 <= 32'h681BA758;
        10'd236 : X0 <= 32'h68068068;
        10'd237 : X0 <= 32'h67F1620E;
        10'd238 : X0 <= 32'h67DC4C46;
        10'd239 : X0 <= 32'h67C73F0A;
        10'd240 : X0 <= 32'h67B23A54;
        10'd241 : X0 <= 32'h679D3E21;
        10'd242 : X0 <= 32'h67884A6A;
        10'd243 : X0 <= 32'h67735F2B;
        10'd244 : X0 <= 32'h675E7C5E;
        10'd245 : X0 <= 32'h6749A1FE;
        10'd246 : X0 <= 32'h6734D006;
        10'd247 : X0 <= 32'h67200672;
        10'd248 : X0 <= 32'h670B453C;
        10'd249 : X0 <= 32'h66F68C5E;
        10'd250 : X0 <= 32'h66E1DBD5;
        10'd251 : X0 <= 32'h66CD339A;
        10'd252 : X0 <= 32'h66B893A9;
        10'd253 : X0 <= 32'h66A3FBFE;
        10'd254 : X0 <= 32'h668F6C92;
        10'd255 : X0 <= 32'h667AE561;
        10'd256 : X0 <= 32'h66666666;
        10'd257 : X0 <= 32'h6651EF9D;
        10'd258 : X0 <= 32'h663D8100;
        10'd259 : X0 <= 32'h66291A8A;
        10'd260 : X0 <= 32'h6614BC36;
        10'd261 : X0 <= 32'h66006600;
        10'd262 : X0 <= 32'h65EC17E3;
        10'd263 : X0 <= 32'h65D7D1DA;
        10'd264 : X0 <= 32'h65C393E0;
        10'd265 : X0 <= 32'h65AF5DF1;
        10'd266 : X0 <= 32'h659B3006;
        10'd267 : X0 <= 32'h65870A1D;
        10'd268 : X0 <= 32'h6572EC30;
        10'd269 : X0 <= 32'h655ED639;
        10'd270 : X0 <= 32'h654AC836;
        10'd271 : X0 <= 32'h6536C220;
        10'd272 : X0 <= 32'h6522C3F3;
        10'd273 : X0 <= 32'h650ECDAB;
        10'd274 : X0 <= 32'h64FADF43;
        10'd275 : X0 <= 32'h64E6F8B5;
        10'd276 : X0 <= 32'h64D319FE;
        10'd277 : X0 <= 32'h64BF4319;
        10'd278 : X0 <= 32'h64AB7402;
        10'd279 : X0 <= 32'h6497ACB2;
        10'd280 : X0 <= 32'h6483ED27;
        10'd281 : X0 <= 32'h6470355C;
        10'd282 : X0 <= 32'h645C854B;
        10'd283 : X0 <= 32'h6448DCF1;
        10'd284 : X0 <= 32'h64353C48;
        10'd285 : X0 <= 32'h6421A34D;
        10'd286 : X0 <= 32'h640E11FB;
        10'd287 : X0 <= 32'h63FA884D;
        10'd288 : X0 <= 32'h63E7063E;
        10'd289 : X0 <= 32'h63D38BCC;
        10'd290 : X0 <= 32'h63C018F0;
        10'd291 : X0 <= 32'h63ACADA7;
        10'd292 : X0 <= 32'h639949EC;
        10'd293 : X0 <= 32'h6385EDBA;
        10'd294 : X0 <= 32'h6372990E;
        10'd295 : X0 <= 32'h635F4BE3;
        10'd296 : X0 <= 32'h634C0635;
        10'd297 : X0 <= 32'h6338C7FE;
        10'd298 : X0 <= 32'h6325913C;
        10'd299 : X0 <= 32'h631261E9;
        10'd300 : X0 <= 32'h62FF3A02;
        10'd301 : X0 <= 32'h62EC1981;
        10'd302 : X0 <= 32'h62D90063;
        10'd303 : X0 <= 32'h62C5EEA3;
        10'd304 : X0 <= 32'h62B2E43E;
        10'd305 : X0 <= 32'h629FE12E;
        10'd306 : X0 <= 32'h628CE570;
        10'd307 : X0 <= 32'h6279F0FF;
        10'd308 : X0 <= 32'h626703D8;
        10'd309 : X0 <= 32'h62541DF6;
        10'd310 : X0 <= 32'h62413F54;
        10'd311 : X0 <= 32'h622E67EF;
        10'd312 : X0 <= 32'h621B97C3;
        10'd313 : X0 <= 32'h6208CECB;
        10'd314 : X0 <= 32'h61F60D03;
        10'd315 : X0 <= 32'h61E35267;
        10'd316 : X0 <= 32'h61D09EF3;
        10'd317 : X0 <= 32'h61BDF2A3;
        10'd318 : X0 <= 32'h61AB4D73;
        10'd319 : X0 <= 32'h6198AF5E;
        10'd320 : X0 <= 32'h61861862;
        10'd321 : X0 <= 32'h61738878;
        10'd322 : X0 <= 32'h6160FF9F;
        10'd323 : X0 <= 32'h614E7DD0;
        10'd324 : X0 <= 32'h613C030A;
        10'd325 : X0 <= 32'h61298F47;
        10'd326 : X0 <= 32'h61172283;
        10'd327 : X0 <= 32'h6104BCBB;
        10'd328 : X0 <= 32'h60F25DEB;
        10'd329 : X0 <= 32'h60E0060E;
        10'd330 : X0 <= 32'h60CDB521;
        10'd331 : X0 <= 32'h60BB6B20;
        10'd332 : X0 <= 32'h60A92806;
        10'd333 : X0 <= 32'h6096EBD0;
        10'd334 : X0 <= 32'h6084B67B;
        10'd335 : X0 <= 32'h60728802;
        10'd336 : X0 <= 32'h60606060;
        10'd337 : X0 <= 32'h604E3F94;
        10'd338 : X0 <= 32'h603C2597;
        10'd339 : X0 <= 32'h602A1268;
        10'd340 : X0 <= 32'h60180602;
        10'd341 : X0 <= 32'h60060060;
        10'd342 : X0 <= 32'h5FF40180;
        10'd343 : X0 <= 32'h5FE2095D;
        10'd344 : X0 <= 32'h5FD017F4;
        10'd345 : X0 <= 32'h5FBE2D41;
        10'd346 : X0 <= 32'h5FAC4940;
        10'd347 : X0 <= 32'h5F9A6BED;
        10'd348 : X0 <= 32'h5F889545;
        10'd349 : X0 <= 32'h5F76C544;
        10'd350 : X0 <= 32'h5F64FBE7;
        10'd351 : X0 <= 32'h5F533928;
        10'd352 : X0 <= 32'h5F417D06;
        10'd353 : X0 <= 32'h5F2FC77C;
        10'd354 : X0 <= 32'h5F1E1886;
        10'd355 : X0 <= 32'h5F0C7021;
        10'd356 : X0 <= 32'h5EFACE49;
        10'd357 : X0 <= 32'h5EE932FA;
        10'd358 : X0 <= 32'h5ED79E32;
        10'd359 : X0 <= 32'h5EC60FEB;
        10'd360 : X0 <= 32'h5EB48824;
        10'd361 : X0 <= 32'h5EA306D7;
        10'd362 : X0 <= 32'h5E918C01;
        10'd363 : X0 <= 32'h5E8017A0;
        10'd364 : X0 <= 32'h5E6EA9AF;
        10'd365 : X0 <= 32'h5E5D422A;
        10'd366 : X0 <= 32'h5E4BE10F;
        10'd367 : X0 <= 32'h5E3A8659;
        10'd368 : X0 <= 32'h5E293206;
        10'd369 : X0 <= 32'h5E17E411;
        10'd370 : X0 <= 32'h5E069C77;
        10'd371 : X0 <= 32'h5DF55B35;
        10'd372 : X0 <= 32'h5DE42046;
        10'd373 : X0 <= 32'h5DD2EBA9;
        10'd374 : X0 <= 32'h5DC1BD58;
        10'd375 : X0 <= 32'h5DB09551;
        10'd376 : X0 <= 32'h5D9F7391;
        10'd377 : X0 <= 32'h5D8E5813;
        10'd378 : X0 <= 32'h5D7D42D5;
        10'd379 : X0 <= 32'h5D6C33D2;
        10'd380 : X0 <= 32'h5D5B2B08;
        10'd381 : X0 <= 32'h5D4A2873;
        10'd382 : X0 <= 32'h5D392C10;
        10'd383 : X0 <= 32'h5D2835DB;
        10'd384 : X0 <= 32'h5D1745D1;
        10'd385 : X0 <= 32'h5D065BEF;
        10'd386 : X0 <= 32'h5CF57831;
        10'd387 : X0 <= 32'h5CE49A94;
        10'd388 : X0 <= 32'h5CD3C315;
        10'd389 : X0 <= 32'h5CC2F1B0;
        10'd390 : X0 <= 32'h5CB22662;
        10'd391 : X0 <= 32'h5CA16127;
        10'd392 : X0 <= 32'h5C90A1FD;
        10'd393 : X0 <= 32'h5C7FE8E0;
        10'd394 : X0 <= 32'h5C6F35CD;
        10'd395 : X0 <= 32'h5C5E88C0;
        10'd396 : X0 <= 32'h5C4DE1B6;
        10'd397 : X0 <= 32'h5C3D40AD;
        10'd398 : X0 <= 32'h5C2CA5A0;
        10'd399 : X0 <= 32'h5C1C108D;
        10'd400 : X0 <= 32'h5C0B8170;
        10'd401 : X0 <= 32'h5BFAF846;
        10'd402 : X0 <= 32'h5BEA750D;
        10'd403 : X0 <= 32'h5BD9F7BF;
        10'd404 : X0 <= 32'h5BC9805C;
        10'd405 : X0 <= 32'h5BB90EDE;
        10'd406 : X0 <= 32'h5BA8A344;
        10'd407 : X0 <= 32'h5B983D8A;
        10'd408 : X0 <= 32'h5B87DDAD;
        10'd409 : X0 <= 32'h5B7783AA;
        10'd410 : X0 <= 32'h5B672F7D;
        10'd411 : X0 <= 32'h5B56E123;
        10'd412 : X0 <= 32'h5B46989A;
        10'd413 : X0 <= 32'h5B3655DE;
        10'd414 : X0 <= 32'h5B2618EC;
        10'd415 : X0 <= 32'h5B15E1C2;
        10'd416 : X0 <= 32'h5B05B05B;
        10'd417 : X0 <= 32'h5AF584B5;
        10'd418 : X0 <= 32'h5AE55ECD;
        10'd419 : X0 <= 32'h5AD53EA0;
        10'd420 : X0 <= 32'h5AC5242B;
        10'd421 : X0 <= 32'h5AB50F6A;
        10'd422 : X0 <= 32'h5AA5005B;
        10'd423 : X0 <= 32'h5A94F6FA;
        10'd424 : X0 <= 32'h5A84F345;
        10'd425 : X0 <= 32'h5A74F539;
        10'd426 : X0 <= 32'h5A64FCD2;
        10'd427 : X0 <= 32'h5A550A0E;
        10'd428 : X0 <= 32'h5A451CEA;
        10'd429 : X0 <= 32'h5A353562;
        10'd430 : X0 <= 32'h5A255375;
        10'd431 : X0 <= 32'h5A15771D;
        10'd432 : X0 <= 32'h5A05A05A;
        10'd433 : X0 <= 32'h59F5CF28;
        10'd434 : X0 <= 32'h59E60383;
        10'd435 : X0 <= 32'h59D63D69;
        10'd436 : X0 <= 32'h59C67CD8;
        10'd437 : X0 <= 32'h59B6C1CC;
        10'd438 : X0 <= 32'h59A70C42;
        10'd439 : X0 <= 32'h59975C37;
        10'd440 : X0 <= 32'h5987B1A9;
        10'd441 : X0 <= 32'h59780C95;
        10'd442 : X0 <= 32'h59686CF7;
        10'd443 : X0 <= 32'h5958D2CE;
        10'd444 : X0 <= 32'h59493E15;
        10'd445 : X0 <= 32'h5939AECA;
        10'd446 : X0 <= 32'h592A24EB;
        10'd447 : X0 <= 32'h591AA075;
        10'd448 : X0 <= 32'h590B2164;
        10'd449 : X0 <= 32'h58FBA7B6;
        10'd450 : X0 <= 32'h58EC3369;
        10'd451 : X0 <= 32'h58DCC478;
        10'd452 : X0 <= 32'h58CD5AE2;
        10'd453 : X0 <= 32'h58BDF6A4;
        10'd454 : X0 <= 32'h58AE97BB;
        10'd455 : X0 <= 32'h589F3E24;
        10'd456 : X0 <= 32'h588FE9DC;
        10'd457 : X0 <= 32'h58809AE1;
        10'd458 : X0 <= 32'h58715130;
        10'd459 : X0 <= 32'h58620CC6;
        10'd460 : X0 <= 32'h5852CDA1;
        10'd461 : X0 <= 32'h584393BD;
        10'd462 : X0 <= 32'h58345F18;
        10'd463 : X0 <= 32'h58252FB0;
        10'd464 : X0 <= 32'h58160581;
        10'd465 : X0 <= 32'h5806E08A;
        10'd466 : X0 <= 32'h57F7C0C6;
        10'd467 : X0 <= 32'h57E8A634;
        10'd468 : X0 <= 32'h57D990D1;
        10'd469 : X0 <= 32'h57CA809A;
        10'd470 : X0 <= 32'h57BB758C;
        10'd471 : X0 <= 32'h57AC6FA6;
        10'd472 : X0 <= 32'h579D6EE3;
        10'd473 : X0 <= 32'h578E7343;
        10'd474 : X0 <= 32'h577F7CC1;
        10'd475 : X0 <= 32'h57708B5B;
        10'd476 : X0 <= 32'h57619F10;
        10'd477 : X0 <= 32'h5752B7DB;
        10'd478 : X0 <= 32'h5743D5BB;
        10'd479 : X0 <= 32'h5734F8AD;
        10'd480 : X0 <= 32'h572620AE;
        10'd481 : X0 <= 32'h57174DBC;
        10'd482 : X0 <= 32'h57087FD4;
        10'd483 : X0 <= 32'h56F9B6F4;
        10'd484 : X0 <= 32'h56EAF319;
        10'd485 : X0 <= 32'h56DC3440;
        10'd486 : X0 <= 32'h56CD7A68;
        10'd487 : X0 <= 32'h56BEC58C;
        10'd488 : X0 <= 32'h56B015AC;
        10'd489 : X0 <= 32'h56A16AC4;
        10'd490 : X0 <= 32'h5692C4D2;
        10'd491 : X0 <= 32'h568423D3;
        10'd492 : X0 <= 32'h567587C5;
        10'd493 : X0 <= 32'h5666F0A5;
        10'd494 : X0 <= 32'h56585E71;
        10'd495 : X0 <= 32'h5649D126;
        10'd496 : X0 <= 32'h563B48C2;
        10'd497 : X0 <= 32'h562CC542;
        10'd498 : X0 <= 32'h561E46A5;
        10'd499 : X0 <= 32'h560FCCE7;
        10'd500 : X0 <= 32'h56015805;
        10'd501 : X0 <= 32'h55F2E7FF;
        10'd502 : X0 <= 32'h55E47CD0;
        10'd503 : X0 <= 32'h55D61677;
        10'd504 : X0 <= 32'h55C7B4F1;
        10'd505 : X0 <= 32'h55B9583C;
        10'd506 : X0 <= 32'h55AB0056;
        10'd507 : X0 <= 32'h559CAD3B;
        10'd508 : X0 <= 32'h558E5EEA;
        10'd509 : X0 <= 32'h55801560;
        10'd510 : X0 <= 32'h5571D09B;
        10'd511 : X0 <= 32'h55639098;
        10'd512 : X0 <= 32'h55555555;
        10'd513 : X0 <= 32'h55471ED0;
        10'd514 : X0 <= 32'h5538ED06;
        10'd515 : X0 <= 32'h552ABFF5;
        10'd516 : X0 <= 32'h551C979B;
        10'd517 : X0 <= 32'h550E73F5;
        10'd518 : X0 <= 32'h55005500;
        10'd519 : X0 <= 32'h54F23ABB;
        10'd520 : X0 <= 32'h54E42524;
        10'd521 : X0 <= 32'h54D61437;
        10'd522 : X0 <= 32'h54C807F3;
        10'd523 : X0 <= 32'h54BA0055;
        10'd524 : X0 <= 32'h54ABFD5B;
        10'd525 : X0 <= 32'h549DFF02;
        10'd526 : X0 <= 32'h54900549;
        10'd527 : X0 <= 32'h5482102D;
        10'd528 : X0 <= 32'h54741FAC;
        10'd529 : X0 <= 32'h546633C3;
        10'd530 : X0 <= 32'h54584C70;
        10'd531 : X0 <= 32'h544A69B1;
        10'd532 : X0 <= 32'h543C8B84;
        10'd533 : X0 <= 32'h542EB1E7;
        10'd534 : X0 <= 32'h5420DCD6;
        10'd535 : X0 <= 32'h54130C51;
        10'd536 : X0 <= 32'h54054054;
        10'd537 : X0 <= 32'h53F778DE;
        10'd538 : X0 <= 32'h53E9B5EC;
        10'd539 : X0 <= 32'h53DBF77C;
        10'd540 : X0 <= 32'h53CE3D8B;
        10'd541 : X0 <= 32'h53C08819;
        10'd542 : X0 <= 32'h53B2D722;
        10'd543 : X0 <= 32'h53A52AA4;
        10'd544 : X0 <= 32'h5397829D;
        10'd545 : X0 <= 32'h5389DF0B;
        10'd546 : X0 <= 32'h537C3FEB;
        10'd547 : X0 <= 32'h536EA53C;
        10'd548 : X0 <= 32'h53610EFB;
        10'd549 : X0 <= 32'h53537D27;
        10'd550 : X0 <= 32'h5345EFBC;
        10'd551 : X0 <= 32'h533866BA;
        10'd552 : X0 <= 32'h532AE21D;
        10'd553 : X0 <= 32'h531D61E3;
        10'd554 : X0 <= 32'h530FE60B;
        10'd555 : X0 <= 32'h53026E92;
        10'd556 : X0 <= 32'h52F4FB77;
        10'd557 : X0 <= 32'h52E78CB6;
        10'd558 : X0 <= 32'h52DA224E;
        10'd559 : X0 <= 32'h52CCBC3D;
        10'd560 : X0 <= 32'h52BF5A81;
        10'd561 : X0 <= 32'h52B1FD18;
        10'd562 : X0 <= 32'h52A4A3FF;
        10'd563 : X0 <= 32'h52974F34;
        10'd564 : X0 <= 32'h5289FEB6;
        10'd565 : X0 <= 32'h527CB282;
        10'd566 : X0 <= 32'h526F6A96;
        10'd567 : X0 <= 32'h526226F0;
        10'd568 : X0 <= 32'h5254E78F;
        10'd569 : X0 <= 32'h5247AC6F;
        10'd570 : X0 <= 32'h523A7590;
        10'd571 : X0 <= 32'h522D42EE;
        10'd572 : X0 <= 32'h52201488;
        10'd573 : X0 <= 32'h5212EA5C;
        10'd574 : X0 <= 32'h5205C468;
        10'd575 : X0 <= 32'h51F8A2A9;
        10'd576 : X0 <= 32'h51EB851F;
        10'd577 : X0 <= 32'h51DE6BC6;
        10'd578 : X0 <= 32'h51D1569D;
        10'd579 : X0 <= 32'h51C445A1;
        10'd580 : X0 <= 32'h51B738D1;
        10'd581 : X0 <= 32'h51AA302B;
        10'd582 : X0 <= 32'h519D2BAD;
        10'd583 : X0 <= 32'h51902B55;
        10'd584 : X0 <= 32'h51832F20;
        10'd585 : X0 <= 32'h5176370D;
        10'd586 : X0 <= 32'h5169431A;
        10'd587 : X0 <= 32'h515C5344;
        10'd588 : X0 <= 32'h514F678B;
        10'd589 : X0 <= 32'h51427FEC;
        10'd590 : X0 <= 32'h51359C64;
        10'd591 : X0 <= 32'h5128BCF3;
        10'd592 : X0 <= 32'h511BE196;
        10'd593 : X0 <= 32'h510F0A4A;
        10'd594 : X0 <= 32'h51023710;
        10'd595 : X0 <= 32'h50F567E3;
        10'd596 : X0 <= 32'h50E89CC3;
        10'd597 : X0 <= 32'h50DBD5AD;
        10'd598 : X0 <= 32'h50CF12A0;
        10'd599 : X0 <= 32'h50C25399;
        10'd600 : X0 <= 32'h50B59897;
        10'd601 : X0 <= 32'h50A8E198;
        10'd602 : X0 <= 32'h509C2E9A;
        10'd603 : X0 <= 32'h508F7F9B;
        10'd604 : X0 <= 32'h5082D499;
        10'd605 : X0 <= 32'h50762D93;
        10'd606 : X0 <= 32'h50698A86;
        10'd607 : X0 <= 32'h505CEB70;
        10'd608 : X0 <= 32'h50505050;
        10'd609 : X0 <= 32'h5043B924;
        10'd610 : X0 <= 32'h503725EA;
        10'd611 : X0 <= 32'h502A96A0;
        10'd612 : X0 <= 32'h501E0B44;
        10'd613 : X0 <= 32'h501183D5;
        10'd614 : X0 <= 32'h50050050;
        10'd615 : X0 <= 32'h4FF880B4;
        10'd616 : X0 <= 32'h4FEC04FF;
        10'd617 : X0 <= 32'h4FDF8D2F;
        10'd618 : X0 <= 32'h4FD31942;
        10'd619 : X0 <= 32'h4FC6A936;
        10'd620 : X0 <= 32'h4FBA3D0B;
        10'd621 : X0 <= 32'h4FADD4BD;
        10'd622 : X0 <= 32'h4FA1704B;
        10'd623 : X0 <= 32'h4F950FB3;
        10'd624 : X0 <= 32'h4F88B2F4;
        10'd625 : X0 <= 32'h4F7C5A0B;
        10'd626 : X0 <= 32'h4F7004F7;
        10'd627 : X0 <= 32'h4F63B3B6;
        10'd628 : X0 <= 32'h4F576647;
        10'd629 : X0 <= 32'h4F4B1CA7;
        10'd630 : X0 <= 32'h4F3ED6D4;
        10'd631 : X0 <= 32'h4F3294CE;
        10'd632 : X0 <= 32'h4F265692;
        10'd633 : X0 <= 32'h4F1A1C1E;
        10'd634 : X0 <= 32'h4F0DE571;
        10'd635 : X0 <= 32'h4F01B289;
        10'd636 : X0 <= 32'h4EF58365;
        10'd637 : X0 <= 32'h4EE95801;
        10'd638 : X0 <= 32'h4EDD305E;
        10'd639 : X0 <= 32'h4ED10C78;
        10'd640 : X0 <= 32'h4EC4EC4F;
        10'd641 : X0 <= 32'h4EB8CFE0;
        10'd642 : X0 <= 32'h4EACB72A;
        10'd643 : X0 <= 32'h4EA0A22B;
        10'd644 : X0 <= 32'h4E9490E2;
        10'd645 : X0 <= 32'h4E88834C;
        10'd646 : X0 <= 32'h4E7C7969;
        10'd647 : X0 <= 32'h4E707335;
        10'd648 : X0 <= 32'h4E6470B0;
        10'd649 : X0 <= 32'h4E5871D9;
        10'd650 : X0 <= 32'h4E4C76AC;
        10'd651 : X0 <= 32'h4E407F29;
        10'd652 : X0 <= 32'h4E348B4E;
        10'd653 : X0 <= 32'h4E289B19;
        10'd654 : X0 <= 32'h4E1CAE88;
        10'd655 : X0 <= 32'h4E10C59A;
        10'd656 : X0 <= 32'h4E04E04E;
        10'd657 : X0 <= 32'h4DF8FEA1;
        10'd658 : X0 <= 32'h4DED2092;
        10'd659 : X0 <= 32'h4DE1461F;
        10'd660 : X0 <= 32'h4DD56F47;
        10'd661 : X0 <= 32'h4DC99C08;
        10'd662 : X0 <= 32'h4DBDCC60;
        10'd663 : X0 <= 32'h4DB2004E;
        10'd664 : X0 <= 32'h4DA637CF;
        10'd665 : X0 <= 32'h4D9A72E4;
        10'd666 : X0 <= 32'h4D8EB189;
        10'd667 : X0 <= 32'h4D82F3BD;
        10'd668 : X0 <= 32'h4D77397E;
        10'd669 : X0 <= 32'h4D6B82CC;
        10'd670 : X0 <= 32'h4D5FCFA4;
        10'd671 : X0 <= 32'h4D542005;
        10'd672 : X0 <= 32'h4D4873ED;
        10'd673 : X0 <= 32'h4D3CCB5A;
        10'd674 : X0 <= 32'h4D31264B;
        10'd675 : X0 <= 32'h4D2584BF;
        10'd676 : X0 <= 32'h4D19E6B4;
        10'd677 : X0 <= 32'h4D0E4C27;
        10'd678 : X0 <= 32'h4D02B518;
        10'd679 : X0 <= 32'h4CF72186;
        10'd680 : X0 <= 32'h4CEB916D;
        10'd681 : X0 <= 32'h4CE004CE;
        10'd682 : X0 <= 32'h4CD47BA6;
        10'd683 : X0 <= 32'h4CC8F5F4;
        10'd684 : X0 <= 32'h4CBD73B6;
        10'd685 : X0 <= 32'h4CB1F4EA;
        10'd686 : X0 <= 32'h4CA67990;
        10'd687 : X0 <= 32'h4C9B01A5;
        10'd688 : X0 <= 32'h4C8F8D29;
        10'd689 : X0 <= 32'h4C841C19;
        10'd690 : X0 <= 32'h4C78AE73;
        10'd691 : X0 <= 32'h4C6D4438;
        10'd692 : X0 <= 32'h4C61DD64;
        10'd693 : X0 <= 32'h4C5679F6;
        10'd694 : X0 <= 32'h4C4B19EE;
        10'd695 : X0 <= 32'h4C3FBD48;
        10'd696 : X0 <= 32'h4C346405;
        10'd697 : X0 <= 32'h4C290E22;
        10'd698 : X0 <= 32'h4C1DBB9D;
        10'd699 : X0 <= 32'h4C126C76;
        10'd700 : X0 <= 32'h4C0720AB;
        10'd701 : X0 <= 32'h4BFBD83A;
        10'd702 : X0 <= 32'h4BF09322;
        10'd703 : X0 <= 32'h4BE55161;
        10'd704 : X0 <= 32'h4BDA12F7;
        10'd705 : X0 <= 32'h4BCED7E0;
        10'd706 : X0 <= 32'h4BC3A01C;
        10'd707 : X0 <= 32'h4BB86BAA;
        10'd708 : X0 <= 32'h4BAD3A88;
        10'd709 : X0 <= 32'h4BA20CB4;
        10'd710 : X0 <= 32'h4B96E22D;
        10'd711 : X0 <= 32'h4B8BBAF2;
        10'd712 : X0 <= 32'h4B809701;
        10'd713 : X0 <= 32'h4B757659;
        10'd714 : X0 <= 32'h4B6A58F7;
        10'd715 : X0 <= 32'h4B5F3EDC;
        10'd716 : X0 <= 32'h4B542805;
        10'd717 : X0 <= 32'h4B491470;
        10'd718 : X0 <= 32'h4B3E041D;
        10'd719 : X0 <= 32'h4B32F70A;
        10'd720 : X0 <= 32'h4B27ED36;
        10'd721 : X0 <= 32'h4B1CE69F;
        10'd722 : X0 <= 32'h4B11E343;
        10'd723 : X0 <= 32'h4B06E322;
        10'd724 : X0 <= 32'h4AFBE639;
        10'd725 : X0 <= 32'h4AF0EC88;
        10'd726 : X0 <= 32'h4AE5F60D;
        10'd727 : X0 <= 32'h4ADB02C7;
        10'd728 : X0 <= 32'h4AD012B4;
        10'd729 : X0 <= 32'h4AC525D3;
        10'd730 : X0 <= 32'h4ABA3C22;
        10'd731 : X0 <= 32'h4AAF55A0;
        10'd732 : X0 <= 32'h4AA4724C;
        10'd733 : X0 <= 32'h4A999224;
        10'd734 : X0 <= 32'h4A8EB527;
        10'd735 : X0 <= 32'h4A83DB53;
        10'd736 : X0 <= 32'h4A7904A8;
        10'd737 : X0 <= 32'h4A6E3123;
        10'd738 : X0 <= 32'h4A6360C3;
        10'd739 : X0 <= 32'h4A589388;
        10'd740 : X0 <= 32'h4A4DC96F;
        10'd741 : X0 <= 32'h4A430277;
        10'd742 : X0 <= 32'h4A383E9F;
        10'd743 : X0 <= 32'h4A2D7DE6;
        10'd744 : X0 <= 32'h4A22C04A;
        10'd745 : X0 <= 32'h4A1805CA;
        10'd746 : X0 <= 32'h4A0D4E64;
        10'd747 : X0 <= 32'h4A029A17;
        10'd748 : X0 <= 32'h49F7E8E3;
        10'd749 : X0 <= 32'h49ED3AC4;
        10'd750 : X0 <= 32'h49E28FBB;
        10'd751 : X0 <= 32'h49D7E7C5;
        10'd752 : X0 <= 32'h49CD42E2;
        10'd753 : X0 <= 32'h49C2A110;
        10'd754 : X0 <= 32'h49B8024E;
        10'd755 : X0 <= 32'h49AD669A;
        10'd756 : X0 <= 32'h49A2CDF3;
        10'd757 : X0 <= 32'h49983859;
        10'd758 : X0 <= 32'h498DA5C8;
        10'd759 : X0 <= 32'h49831641;
        10'd760 : X0 <= 32'h497889C2;
        10'd761 : X0 <= 32'h496E0049;
        10'd762 : X0 <= 32'h496379D6;
        10'd763 : X0 <= 32'h4958F667;
        10'd764 : X0 <= 32'h494E75FA;
        10'd765 : X0 <= 32'h4943F88F;
        10'd766 : X0 <= 32'h49397E24;
        10'd767 : X0 <= 32'h492F06B8;
        10'd768 : X0 <= 32'h49249249;
        10'd769 : X0 <= 32'h491A20D7;
        10'd770 : X0 <= 32'h490FB25F;
        10'd771 : X0 <= 32'h490546E2;
        10'd772 : X0 <= 32'h48FADE5C;
        10'd773 : X0 <= 32'h48F078CE;
        10'd774 : X0 <= 32'h48E61636;
        10'd775 : X0 <= 32'h48DBB693;
        10'd776 : X0 <= 32'h48D159E2;
        10'd777 : X0 <= 32'h48C70024;
        10'd778 : X0 <= 32'h48BCA957;
        10'd779 : X0 <= 32'h48B2557A;
        10'd780 : X0 <= 32'h48A8048B;
        10'd781 : X0 <= 32'h489DB688;
        10'd782 : X0 <= 32'h48936B72;
        10'd783 : X0 <= 32'h48892347;
        10'd784 : X0 <= 32'h487EDE05;
        10'd785 : X0 <= 32'h48749BAB;
        10'd786 : X0 <= 32'h486A5C37;
        10'd787 : X0 <= 32'h48601FAA;
        10'd788 : X0 <= 32'h4855E601;
        10'd789 : X0 <= 32'h484BAF3B;
        10'd790 : X0 <= 32'h48417B58;
        10'd791 : X0 <= 32'h48374A55;
        10'd792 : X0 <= 32'h482D1C32;
        10'd793 : X0 <= 32'h4822F0ED;
        10'd794 : X0 <= 32'h4818C885;
        10'd795 : X0 <= 32'h480EA2F9;
        10'd796 : X0 <= 32'h48048048;
        10'd797 : X0 <= 32'h47FA6070;
        10'd798 : X0 <= 32'h47F04371;
        10'd799 : X0 <= 32'h47E62949;
        10'd800 : X0 <= 32'h47DC11F7;
        10'd801 : X0 <= 32'h47D1FD7A;
        10'd802 : X0 <= 32'h47C7EBD0;
        10'd803 : X0 <= 32'h47BDDCF8;
        10'd804 : X0 <= 32'h47B3D0F2;
        10'd805 : X0 <= 32'h47A9C7BC;
        10'd806 : X0 <= 32'h479FC154;
        10'd807 : X0 <= 32'h4795BDBA;
        10'd808 : X0 <= 32'h478BBCED;
        10'd809 : X0 <= 32'h4781BEEB;
        10'd810 : X0 <= 32'h4777C3B3;
        10'd811 : X0 <= 32'h476DCB44;
        10'd812 : X0 <= 32'h4763D59D;
        10'd813 : X0 <= 32'h4759E2BC;
        10'd814 : X0 <= 32'h474FF2A1;
        10'd815 : X0 <= 32'h4746054A;
        10'd816 : X0 <= 32'h473C1AB7;
        10'd817 : X0 <= 32'h473232E5;
        10'd818 : X0 <= 32'h47284DD4;
        10'd819 : X0 <= 32'h471E6B83;
        10'd820 : X0 <= 32'h47148BF0;
        10'd821 : X0 <= 32'h470AAF1B;
        10'd822 : X0 <= 32'h4700D502;
        10'd823 : X0 <= 32'h46F6FDA5;
        10'd824 : X0 <= 32'h46ED2901;
        10'd825 : X0 <= 32'h46E35716;
        10'd826 : X0 <= 32'h46D987E3;
        10'd827 : X0 <= 32'h46CFBB67;
        10'd828 : X0 <= 32'h46C5F1A0;
        10'd829 : X0 <= 32'h46BC2A8D;
        10'd830 : X0 <= 32'h46B2662E;
        10'd831 : X0 <= 32'h46A8A481;
        10'd832 : X0 <= 32'h469EE584;
        10'd833 : X0 <= 32'h46952938;
        10'd834 : X0 <= 32'h468B6F9B;
        10'd835 : X0 <= 32'h4681B8AB;
        10'd836 : X0 <= 32'h46780468;
        10'd837 : X0 <= 32'h466E52D0;
        10'd838 : X0 <= 32'h4664A3E2;
        10'd839 : X0 <= 32'h465AF79E;
        10'd840 : X0 <= 32'h46514E02;
        10'd841 : X0 <= 32'h4647A70D;
        10'd842 : X0 <= 32'h463E02BE;
        10'd843 : X0 <= 32'h46346114;
        10'd844 : X0 <= 32'h462AC20E;
        10'd845 : X0 <= 32'h462125AB;
        10'd846 : X0 <= 32'h46178BE9;
        10'd847 : X0 <= 32'h460DF4C8;
        10'd848 : X0 <= 32'h46046046;
        10'd849 : X0 <= 32'h45FACE63;
        10'd850 : X0 <= 32'h45F13F1D;
        10'd851 : X0 <= 32'h45E7B273;
        10'd852 : X0 <= 32'h45DE2864;
        10'd853 : X0 <= 32'h45D4A0F0;
        10'd854 : X0 <= 32'h45CB1C15;
        10'd855 : X0 <= 32'h45C199D1;
        10'd856 : X0 <= 32'h45B81A25;
        10'd857 : X0 <= 32'h45AE9D0F;
        10'd858 : X0 <= 32'h45A5228D;
        10'd859 : X0 <= 32'h459BAA9F;
        10'd860 : X0 <= 32'h45923544;
        10'd861 : X0 <= 32'h4588C27A;
        10'd862 : X0 <= 32'h457F5242;
        10'd863 : X0 <= 32'h4575E498;
        10'd864 : X0 <= 32'h456C797E;
        10'd865 : X0 <= 32'h456310F1;
        10'd866 : X0 <= 32'h4559AAF0;
        10'd867 : X0 <= 32'h4550477B;
        10'd868 : X0 <= 32'h4546E690;
        10'd869 : X0 <= 32'h453D882F;
        10'd870 : X0 <= 32'h45342C55;
        10'd871 : X0 <= 32'h452AD304;
        10'd872 : X0 <= 32'h45217C38;
        10'd873 : X0 <= 32'h451827F2;
        10'd874 : X0 <= 32'h450ED630;
        10'd875 : X0 <= 32'h450586F1;
        10'd876 : X0 <= 32'h44FC3A35;
        10'd877 : X0 <= 32'h44F2EFFA;
        10'd878 : X0 <= 32'h44E9A83E;
        10'd879 : X0 <= 32'h44E06303;
        10'd880 : X0 <= 32'h44D72045;
        10'd881 : X0 <= 32'h44CDE004;
        10'd882 : X0 <= 32'h44C4A240;
        10'd883 : X0 <= 32'h44BB66F7;
        10'd884 : X0 <= 32'h44B22E28;
        10'd885 : X0 <= 32'h44A8F7D2;
        10'd886 : X0 <= 32'h449FC3F4;
        10'd887 : X0 <= 32'h4496928E;
        10'd888 : X0 <= 32'h448D639D;
        10'd889 : X0 <= 32'h44843722;
        10'd890 : X0 <= 32'h447B0D1C;
        10'd891 : X0 <= 32'h4471E588;
        10'd892 : X0 <= 32'h4468C067;
        10'd893 : X0 <= 32'h445F9DB7;
        10'd894 : X0 <= 32'h44567D77;
        10'd895 : X0 <= 32'h444D5FA6;
        10'd896 : X0 <= 32'h44444444;
        10'd897 : X0 <= 32'h443B2B50;
        10'd898 : X0 <= 32'h443214C7;
        10'd899 : X0 <= 32'h442900AA;
        10'd900 : X0 <= 32'h441FEEF8;
        10'd901 : X0 <= 32'h4416DFAF;
        10'd902 : X0 <= 32'h440DD2CF;
        10'd903 : X0 <= 32'h4404C856;
        10'd904 : X0 <= 32'h43FBC044;
        10'd905 : X0 <= 32'h43F2BA98;
        10'd906 : X0 <= 32'h43E9B750;
        10'd907 : X0 <= 32'h43E0B66C;
        10'd908 : X0 <= 32'h43D7B7EB;
        10'd909 : X0 <= 32'h43CEBBCC;
        10'd910 : X0 <= 32'h43C5C20D;
        10'd911 : X0 <= 32'h43BCCAAF;
        10'd912 : X0 <= 32'h43B3D5B0;
        10'd913 : X0 <= 32'h43AAE30E;
        10'd914 : X0 <= 32'h43A1F2CA;
        10'd915 : X0 <= 32'h439904E3;
        10'd916 : X0 <= 32'h43901956;
        10'd917 : X0 <= 32'h43873024;
        10'd918 : X0 <= 32'h437E494B;
        10'd919 : X0 <= 32'h437564CB;
        10'd920 : X0 <= 32'h436C82A2;
        10'd921 : X0 <= 32'h4363A2D0;
        10'd922 : X0 <= 32'h435AC554;
        10'd923 : X0 <= 32'h4351EA2C;
        10'd924 : X0 <= 32'h43491159;
        10'd925 : X0 <= 32'h43403AD8;
        10'd926 : X0 <= 32'h433766AA;
        10'd927 : X0 <= 32'h432E94CC;
        10'd928 : X0 <= 32'h4325C53F;
        10'd929 : X0 <= 32'h431CF801;
        10'd930 : X0 <= 32'h43142D12;
        10'd931 : X0 <= 32'h430B6470;
        10'd932 : X0 <= 32'h43029E1A;
        10'd933 : X0 <= 32'h42F9DA10;
        10'd934 : X0 <= 32'h42F11852;
        10'd935 : X0 <= 32'h42E858DD;
        10'd936 : X0 <= 32'h42DF9BB1;
        10'd937 : X0 <= 32'h42D6E0CD;
        10'd938 : X0 <= 32'h42CE2830;
        10'd939 : X0 <= 32'h42C571DA;
        10'd940 : X0 <= 32'h42BCBDC9;
        10'd941 : X0 <= 32'h42B40BFC;
        10'd942 : X0 <= 32'h42AB5C74;
        10'd943 : X0 <= 32'h42A2AF2E;
        10'd944 : X0 <= 32'h429A042A;
        10'd945 : X0 <= 32'h42915B67;
        10'd946 : X0 <= 32'h4288B4E4;
        10'd947 : X0 <= 32'h428010A0;
        10'd948 : X0 <= 32'h42776E9B;
        10'd949 : X0 <= 32'h426ECED3;
        10'd950 : X0 <= 32'h42663148;
        10'd951 : X0 <= 32'h425D95F8;
        10'd952 : X0 <= 32'h4254FCE4;
        10'd953 : X0 <= 32'h424C660A;
        10'd954 : X0 <= 32'h4243D168;
        10'd955 : X0 <= 32'h423B3EFF;
        10'd956 : X0 <= 32'h4232AECE;
        10'd957 : X0 <= 32'h422A20D3;
        10'd958 : X0 <= 32'h4221950E;
        10'd959 : X0 <= 32'h42190B7D;
        10'd960 : X0 <= 32'h42108421;
        10'd961 : X0 <= 32'h4207FEF8;
        10'd962 : X0 <= 32'h41FF7C01;
        10'd963 : X0 <= 32'h41F6FB3C;
        10'd964 : X0 <= 32'h41EE7CA7;
        10'd965 : X0 <= 32'h41E60042;
        10'd966 : X0 <= 32'h41DD860C;
        10'd967 : X0 <= 32'h41D50E04;
        10'd968 : X0 <= 32'h41CC9829;
        10'd969 : X0 <= 32'h41C4247B;
        10'd970 : X0 <= 32'h41BBB2F8;
        10'd971 : X0 <= 32'h41B343A0;
        10'd972 : X0 <= 32'h41AAD672;
        10'd973 : X0 <= 32'h41A26B6D;
        10'd974 : X0 <= 32'h419A0290;
        10'd975 : X0 <= 32'h41919BDB;
        10'd976 : X0 <= 32'h4189374C;
        10'd977 : X0 <= 32'h4180D4E3;
        10'd978 : X0 <= 32'h4178749F;
        10'd979 : X0 <= 32'h4170167F;
        10'd980 : X0 <= 32'h4167BA82;
        10'd981 : X0 <= 32'h415F60A8;
        10'd982 : X0 <= 32'h415708EF;
        10'd983 : X0 <= 32'h414EB357;
        10'd984 : X0 <= 32'h41465FDF;
        10'd985 : X0 <= 32'h413E0E87;
        10'd986 : X0 <= 32'h4135BF4D;
        10'd987 : X0 <= 32'h412D7230;
        10'd988 : X0 <= 32'h41252730;
        10'd989 : X0 <= 32'h411CDE4D;
        10'd990 : X0 <= 32'h41149784;
        10'd991 : X0 <= 32'h410C52D6;
        10'd992 : X0 <= 32'h41041041;
        10'd993 : X0 <= 32'h40FBCFC5;
        10'd994 : X0 <= 32'h40F39161;
        10'd995 : X0 <= 32'h40EB5514;
        10'd996 : X0 <= 32'h40E31ADE;
        10'd997 : X0 <= 32'h40DAE2BD;
        10'd998 : X0 <= 32'h40D2ACB1;
        10'd999 : X0 <= 32'h40CA78B9;
        10'd1000 : X0 <= 32'h40C246D4;
        10'd1001 : X0 <= 32'h40BA1702;
        10'd1002 : X0 <= 32'h40B1E941;
        10'd1003 : X0 <= 32'h40A9BD92;
        10'd1004 : X0 <= 32'h40A193F2;
        10'd1005 : X0 <= 32'h40996C61;
        10'd1006 : X0 <= 32'h409146DF;
        10'd1007 : X0 <= 32'h4089236B;
        10'd1008 : X0 <= 32'h40810204;
        10'd1009 : X0 <= 32'h4078E2A9;
        10'd1010 : X0 <= 32'h4070C559;
        10'd1011 : X0 <= 32'h4068AA14;
        10'd1012 : X0 <= 32'h406090D9;
        10'd1013 : X0 <= 32'h405879A7;
        10'd1014 : X0 <= 32'h4050647E;
        10'd1015 : X0 <= 32'h4048515C;
        10'd1016 : X0 <= 32'h40404040;
        10'd1017 : X0 <= 32'h4038312B;
        10'd1018 : X0 <= 32'h4030241B;
        10'd1019 : X0 <= 32'h40281910;
        10'd1020 : X0 <= 32'h40201008;
        10'd1021 : X0 <= 32'h40180903;
        10'd1022 : X0 <= 32'h40100401;
        10'd1023 : X0 <= 32'h40080100;
        default : X0 <= 32'hFFFFFFFF;
    endcase
end

endmodule
