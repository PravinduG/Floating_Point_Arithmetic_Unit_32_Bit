`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11/27/2025 09:45:09 PM
// Design Name: 
// Module Name: reciprocal_lut
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module reciprocal_lut(
			 input logic  [9:0]														lut_idx
			,output logic [31:0]													X0

    );
		
		always_comb begin
  case(lut_idx)
    10'd0 : X0 <= 32'hFFFFFFFF;
    10'd1 : X0 <= 32'hFFC00FFC;
    10'd2 : X0 <= 32'hFF803FE0;
    10'd3 : X0 <= 32'hFF408F94;
    10'd4 : X0 <= 32'hFF00FF01;
    10'd5 : X0 <= 32'hFEC18E0E;
    10'd6 : X0 <= 32'hFE823CA5;
    10'd7 : X0 <= 32'hFE430AAD;
    10'd8 : X0 <= 32'hFE03F810;
    10'd9 : X0 <= 32'hFDC504B5;
    10'd10 : X0 <= 32'hFD863087;
    10'd11 : X0 <= 32'hFD477B6D;
    10'd12 : X0 <= 32'hFD08E550;
    10'd13 : X0 <= 32'hFCCA6E1A;
    10'd14 : X0 <= 32'hFC8C15B4;
    10'd15 : X0 <= 32'hFC4DDC07;
    10'd16 : X0 <= 32'hFC0FC0FC;
    10'd17 : X0 <= 32'hFBD1C47D;
    10'd18 : X0 <= 32'hFB93E673;
    10'd19 : X0 <= 32'hFB5626C8;
    10'd20 : X0 <= 32'hFB188565;
    10'd21 : X0 <= 32'hFADB0234;
    10'd22 : X0 <= 32'hFA9D9D20;
    10'd23 : X0 <= 32'hFA605611;
    10'd24 : X0 <= 32'hFA232CF2;
    10'd25 : X0 <= 32'hF9E621AE;
    10'd26 : X0 <= 32'hF9A9342D;
    10'd27 : X0 <= 32'hF96C645B;
    10'd28 : X0 <= 32'hF92FB221;
    10'd29 : X0 <= 32'hF8F31D6B;
    10'd30 : X0 <= 32'hF8B6A622;
    10'd31 : X0 <= 32'hF87A4C32;
    10'd32 : X0 <= 32'hF83E0F84;
    10'd33 : X0 <= 32'hF801F004;
    10'd34 : X0 <= 32'hF7C5ED9C;
    10'd35 : X0 <= 32'hF78A0838;
    10'd36 : X0 <= 32'hF74E3FC2;
    10'd37 : X0 <= 32'hF7129426;
    10'd38 : X0 <= 32'hF6D7054E;
    10'd39 : X0 <= 32'hF69B9325;
    10'd40 : X0 <= 32'hF6603D98;
    10'd41 : X0 <= 32'hF6250491;
    10'd42 : X0 <= 32'hF5E9E7FC;
    10'd43 : X0 <= 32'hF5AEE7C4;
    10'd44 : X0 <= 32'hF57403D6;
    10'd45 : X0 <= 32'hF5393C1C;
    10'd46 : X0 <= 32'hF4FE9082;
    10'd47 : X0 <= 32'hF4C400F5;
    10'd48 : X0 <= 32'hF4898D60;
    10'd49 : X0 <= 32'hF44F35AE;
    10'd50 : X0 <= 32'hF414F9CD;
    10'd51 : X0 <= 32'hF3DAD9A9;
    10'd52 : X0 <= 32'hF3A0D52D;
    10'd53 : X0 <= 32'hF366EC45;
    10'd54 : X0 <= 32'hF32D1EDF;
    10'd55 : X0 <= 32'hF2F36CE7;
    10'd56 : X0 <= 32'hF2B9D648;
    10'd57 : X0 <= 32'hF2805AF0;
    10'd58 : X0 <= 32'hF246FACB;
    10'd59 : X0 <= 32'hF20DB5C7;
    10'd60 : X0 <= 32'hF1D48BCF;
    10'd61 : X0 <= 32'hF19B7CD1;
    10'd62 : X0 <= 32'hF16288B9;
    10'd63 : X0 <= 32'hF129AF75;
    10'd64 : X0 <= 32'hF0F0F0F1;
    10'd65 : X0 <= 32'hF0B84D1B;
    10'd66 : X0 <= 32'hF07FC3E0;
    10'd67 : X0 <= 32'hF047552D;
    10'd68 : X0 <= 32'hF00F00F0;
    10'd69 : X0 <= 32'hEFD6C716;
    10'd70 : X0 <= 32'hEF9EA78C;
    10'd71 : X0 <= 32'hEF66A240;
    10'd72 : X0 <= 32'hEF2EB720;
    10'd73 : X0 <= 32'hEEF6E619;
    10'd74 : X0 <= 32'hEEBF2F19;
    10'd75 : X0 <= 32'hEE87920E;
    10'd76 : X0 <= 32'hEE500EE5;
    10'd77 : X0 <= 32'hEE18A58D;
    10'd78 : X0 <= 32'hEDE155F4;
    10'd79 : X0 <= 32'hEDAA2007;
    10'd80 : X0 <= 32'hED7303B6;
    10'd81 : X0 <= 32'hED3C00ED;
    10'd82 : X0 <= 32'hED05179C;
    10'd83 : X0 <= 32'hECCE47B0;
    10'd84 : X0 <= 32'hEC979119;
    10'd85 : X0 <= 32'hEC60F3C4;
    10'd86 : X0 <= 32'hEC2A6FA0;
    10'd87 : X0 <= 32'hEBF4049C;
    10'd88 : X0 <= 32'hEBBDB2A6;
    10'd89 : X0 <= 32'hEB8779AD;
    10'd90 : X0 <= 32'hEB51599F;
    10'd91 : X0 <= 32'hEB1B526D;
    10'd92 : X0 <= 32'hEAE56404;
    10'd93 : X0 <= 32'hEAAF8E53;
    10'd94 : X0 <= 32'hEA79D14A;
    10'd95 : X0 <= 32'hEA442CD7;
    10'd96 : X0 <= 32'hEA0EA0EA;
    10'd97 : X0 <= 32'hE9D92D72;
    10'd98 : X0 <= 32'hE9A3D25E;
    10'd99 : X0 <= 32'hE96E8F9E;
    10'd100 : X0 <= 32'hE9396520;
    10'd101 : X0 <= 32'hE90452D5;
    10'd102 : X0 <= 32'hE8CF58AB;
    10'd103 : X0 <= 32'hE89A7693;
    10'd104 : X0 <= 32'hE865AC7B;
    10'd105 : X0 <= 32'hE830FA55;
    10'd106 : X0 <= 32'hE7FC600E;
    10'd107 : X0 <= 32'hE7C7DD98;
    10'd108 : X0 <= 32'hE79372E2;
    10'd109 : X0 <= 32'hE75F1FDC;
    10'd110 : X0 <= 32'hE72AE475;
    10'd111 : X0 <= 32'hE6F6C09F;
    10'd112 : X0 <= 32'hE6C2B448;
    10'd113 : X0 <= 32'hE68EBF61;
    10'd114 : X0 <= 32'hE65AE1DB;
    10'd115 : X0 <= 32'hE6271BA5;
    10'd116 : X0 <= 32'hE5F36CB0;
    10'd117 : X0 <= 32'hE5BFD4EC;
    10'd118 : X0 <= 32'hE58C544A;
    10'd119 : X0 <= 32'hE558EAB9;
    10'd120 : X0 <= 32'hE525982B;
    10'd121 : X0 <= 32'hE4F25C90;
    10'd122 : X0 <= 32'hE4BF37D9;
    10'd123 : X0 <= 32'hE48C29F6;
    10'd124 : X0 <= 32'hE45932D8;
    10'd125 : X0 <= 32'hE4265270;
    10'd126 : X0 <= 32'hE3F388AF;
    10'd127 : X0 <= 32'hE3C0D585;
    10'd128 : X0 <= 32'hE38E38E4;
    10'd129 : X0 <= 32'hE35BB2BC;
    10'd130 : X0 <= 32'hE32942FF;
    10'd131 : X0 <= 32'hE2F6E99D;
    10'd132 : X0 <= 32'hE2C4A688;
    10'd133 : X0 <= 32'hE29279B2;
    10'd134 : X0 <= 32'hE260630A;
    10'd135 : X0 <= 32'hE22E6283;
    10'd136 : X0 <= 32'hE1FC780E;
    10'd137 : X0 <= 32'hE1CAA39C;
    10'd138 : X0 <= 32'hE198E51F;
    10'd139 : X0 <= 32'hE1673C88;
    10'd140 : X0 <= 32'hE135A9C9;
    10'd141 : X0 <= 32'hE1042CD4;
    10'd142 : X0 <= 32'hE0D2C599;
    10'd143 : X0 <= 32'hE0A1740B;
    10'd144 : X0 <= 32'hE070381C;
    10'd145 : X0 <= 32'hE03F11BD;
    10'd146 : X0 <= 32'hE00E00E0;
    10'd147 : X0 <= 32'hDFDD0577;
    10'd148 : X0 <= 32'hDFAC1F74;
    10'd149 : X0 <= 32'hDF7B4EC9;
    10'd150 : X0 <= 32'hDF4A9368;
    10'd151 : X0 <= 32'hDF19ED43;
    10'd152 : X0 <= 32'hDEE95C4D;
    10'd153 : X0 <= 32'hDEB8E076;
    10'd154 : X0 <= 32'hDE8879B3;
    10'd155 : X0 <= 32'hDE5827F4;
    10'd156 : X0 <= 32'hDE27EB2C;
    10'd157 : X0 <= 32'hDDF7C34E;
    10'd158 : X0 <= 32'hDDC7B04C;
    10'd159 : X0 <= 32'hDD97B219;
    10'd160 : X0 <= 32'hDD67C8A6;
    10'd161 : X0 <= 32'hDD37F3E7;
    10'd162 : X0 <= 32'hDD0833CE;
    10'd163 : X0 <= 32'hDCD8884E;
    10'd164 : X0 <= 32'hDCA8F159;
    10'd165 : X0 <= 32'hDC796EE2;
    10'd166 : X0 <= 32'hDC4A00DC;
    10'd167 : X0 <= 32'hDC1AA73A;
    10'd168 : X0 <= 32'hDBEB61EF;
    10'd169 : X0 <= 32'hDBBC30ED;
    10'd170 : X0 <= 32'hDB8D1427;
    10'd171 : X0 <= 32'hDB5E0B91;
    10'd172 : X0 <= 32'hDB2F171E;
    10'd173 : X0 <= 32'hDB0036C0;
    10'd174 : X0 <= 32'hDAD16A6B;
    10'd175 : X0 <= 32'hDAA2B212;
    10'd176 : X0 <= 32'hDA740DA7;
    10'd177 : X0 <= 32'hDA457D1F;
    10'd178 : X0 <= 32'hDA17006D;
    10'd179 : X0 <= 32'hD9E89784;
    10'd180 : X0 <= 32'hD9BA4257;
    10'd181 : X0 <= 32'hD98C00DA;
    10'd182 : X0 <= 32'hD95DD300;
    10'd183 : X0 <= 32'hD92FB8BC;
    10'd184 : X0 <= 32'hD901B203;
    10'd185 : X0 <= 32'hD8D3BEC8;
    10'd186 : X0 <= 32'hD8A5DEFF;
    10'd187 : X0 <= 32'hD878129A;
    10'd188 : X0 <= 32'hD84A598F;
    10'd189 : X0 <= 32'hD81CB3D0;
    10'd190 : X0 <= 32'hD7EF2151;
    10'd191 : X0 <= 32'hD7C1A207;
    10'd192 : X0 <= 32'hD79435E5;
    10'd193 : X0 <= 32'hD766DCDF;
    10'd194 : X0 <= 32'hD73996E9;
    10'd195 : X0 <= 32'hD70C63F7;
    10'd196 : X0 <= 32'hD6DF43FD;
    10'd197 : X0 <= 32'hD6B236EF;
    10'd198 : X0 <= 32'hD6853CC1;
    10'd199 : X0 <= 32'hD6585567;
    10'd200 : X0 <= 32'hD62B80D6;
    10'd201 : X0 <= 32'hD5FEBF02;
    10'd202 : X0 <= 32'hD5D20FDF;
    10'd203 : X0 <= 32'hD5A57361;
    10'd204 : X0 <= 32'hD578E97C;
    10'd205 : X0 <= 32'hD54C7226;
    10'd206 : X0 <= 32'hD5200D52;
    10'd207 : X0 <= 32'hD4F3BAF5;
    10'd208 : X0 <= 32'hD4C77B03;
    10'd209 : X0 <= 32'hD49B4D72;
    10'd210 : X0 <= 32'hD46F3234;
    10'd211 : X0 <= 32'hD4432940;
    10'd212 : X0 <= 32'hD417328A;
    10'd213 : X0 <= 32'hD3EB4E05;
    10'd214 : X0 <= 32'hD3BF7BA8;
    10'd215 : X0 <= 32'hD393BB67;
    10'd216 : X0 <= 32'hD3680D37;
    10'd217 : X0 <= 32'hD33C710B;
    10'd218 : X0 <= 32'hD310E6DA;
    10'd219 : X0 <= 32'hD2E56E99;
    10'd220 : X0 <= 32'hD2BA083B;
    10'd221 : X0 <= 32'hD28EB3B7;
    10'd222 : X0 <= 32'hD2637100;
    10'd223 : X0 <= 32'hD238400D;
    10'd224 : X0 <= 32'hD20D20D2;
    10'd225 : X0 <= 32'hD1E21344;
    10'd226 : X0 <= 32'hD1B71759;
    10'd227 : X0 <= 32'hD18C2D05;
    10'd228 : X0 <= 32'hD161543E;
    10'd229 : X0 <= 32'hD1368CF9;
    10'd230 : X0 <= 32'hD10BD72C;
    10'd231 : X0 <= 32'hD0E132CB;
    10'd232 : X0 <= 32'hD0B69FCC;
    10'd233 : X0 <= 32'hD08C1E24;
    10'd234 : X0 <= 32'hD061ADC9;
    10'd235 : X0 <= 32'hD0374EB1;
    10'd236 : X0 <= 32'hD00D00D0;
    10'd237 : X0 <= 32'hCFE2C41C;
    10'd238 : X0 <= 32'hCFB8988C;
    10'd239 : X0 <= 32'hCF8E7E13;
    10'd240 : X0 <= 32'hCF6474A9;
    10'd241 : X0 <= 32'hCF3A7C42;
    10'd242 : X0 <= 32'hCF1094D4;
    10'd243 : X0 <= 32'hCEE6BE55;
    10'd244 : X0 <= 32'hCEBCF8BB;
    10'd245 : X0 <= 32'hCE9343FC;
    10'd246 : X0 <= 32'hCE69A00D;
    10'd247 : X0 <= 32'hCE400CE4;
    10'd248 : X0 <= 32'hCE168A77;
    10'd249 : X0 <= 32'hCDED18BC;
    10'd250 : X0 <= 32'hCDC3B7A9;
    10'd251 : X0 <= 32'hCD9A6734;
    10'd252 : X0 <= 32'hCD712753;
    10'd253 : X0 <= 32'hCD47F7FB;
    10'd254 : X0 <= 32'hCD1ED924;
    10'd255 : X0 <= 32'hCCF5CAC2;
    10'd256 : X0 <= 32'hCCCCCCCD;
    10'd257 : X0 <= 32'hCCA3DF3A;
    10'd258 : X0 <= 32'hCC7B01FF;
    10'd259 : X0 <= 32'hCC523513;
    10'd260 : X0 <= 32'hCC29786C;
    10'd261 : X0 <= 32'hCC00CC01;
    10'd262 : X0 <= 32'hCBD82FC7;
    10'd263 : X0 <= 32'hCBAFA3B4;
    10'd264 : X0 <= 32'hCB8727C0;
    10'd265 : X0 <= 32'hCB5EBBE1;
    10'd266 : X0 <= 32'hCB36600D;
    10'd267 : X0 <= 32'hCB0E143A;
    10'd268 : X0 <= 32'hCAE5D85F;
    10'd269 : X0 <= 32'hCABDAC73;
    10'd270 : X0 <= 32'hCA95906C;
    10'd271 : X0 <= 32'hCA6D8440;
    10'd272 : X0 <= 32'hCA4587E7;
    10'd273 : X0 <= 32'hCA1D9B56;
    10'd274 : X0 <= 32'hC9F5BE85;
    10'd275 : X0 <= 32'hC9CDF16B;
    10'd276 : X0 <= 32'hC9A633FD;
    10'd277 : X0 <= 32'hC97E8633;
    10'd278 : X0 <= 32'hC956E803;
    10'd279 : X0 <= 32'hC92F5965;
    10'd280 : X0 <= 32'hC907DA4F;
    10'd281 : X0 <= 32'hC8E06AB7;
    10'd282 : X0 <= 32'hC8B90A96;
    10'd283 : X0 <= 32'hC891B9E1;
    10'd284 : X0 <= 32'hC86A7890;
    10'd285 : X0 <= 32'hC843469A;
    10'd286 : X0 <= 32'hC81C23F5;
    10'd287 : X0 <= 32'hC7F51099;
    10'd288 : X0 <= 32'hC7CE0C7D;
    10'd289 : X0 <= 32'hC7A71797;
    10'd290 : X0 <= 32'hC78031E0;
    10'd291 : X0 <= 32'hC7595B4E;
    10'd292 : X0 <= 32'hC73293D8;
    10'd293 : X0 <= 32'hC70BDB75;
    10'd294 : X0 <= 32'hC6E5321D;
    10'd295 : X0 <= 32'hC6BE97C7;
    10'd296 : X0 <= 32'hC6980C6A;
    10'd297 : X0 <= 32'hC6718FFD;
    10'd298 : X0 <= 32'hC64B2278;
    10'd299 : X0 <= 32'hC624C3D2;
    10'd300 : X0 <= 32'hC5FE7403;
    10'd301 : X0 <= 32'hC5D83302;
    10'd302 : X0 <= 32'hC5B200C6;
    10'd303 : X0 <= 32'hC58BDD46;
    10'd304 : X0 <= 32'hC565C87B;
    10'd305 : X0 <= 32'hC53FC25C;
    10'd306 : X0 <= 32'hC519CAE0;
    10'd307 : X0 <= 32'hC4F3E1FF;
    10'd308 : X0 <= 32'hC4CE07B0;
    10'd309 : X0 <= 32'hC4A83BEB;
    10'd310 : X0 <= 32'hC4827EA8;
    10'd311 : X0 <= 32'hC45CCFDE;
    10'd312 : X0 <= 32'hC4372F85;
    10'd313 : X0 <= 32'hC4119D95;
    10'd314 : X0 <= 32'hC3EC1A05;
    10'd315 : X0 <= 32'hC3C6A4CE;
    10'd316 : X0 <= 32'hC3A13DE6;
    10'd317 : X0 <= 32'hC37BE546;
    10'd318 : X0 <= 32'hC3569AE6;
    10'd319 : X0 <= 32'hC3315EBD;
    10'd320 : X0 <= 32'hC30C30C3;
    10'd321 : X0 <= 32'hC2E710F1;
    10'd322 : X0 <= 32'hC2C1FF3D;
    10'd323 : X0 <= 32'hC29CFBA1;
    10'd324 : X0 <= 32'hC2780614;
    10'd325 : X0 <= 32'hC2531E8E;
    10'd326 : X0 <= 32'hC22E4506;
    10'd327 : X0 <= 32'hC2097976;
    10'd328 : X0 <= 32'hC1E4BBD6;
    10'd329 : X0 <= 32'hC1C00C1C;
    10'd330 : X0 <= 32'hC19B6A42;
    10'd331 : X0 <= 32'hC176D63F;
    10'd332 : X0 <= 32'hC152500C;
    10'd333 : X0 <= 32'hC12DD7A1;
    10'd334 : X0 <= 32'hC1096CF6;
    10'd335 : X0 <= 32'hC0E51003;
    10'd336 : X0 <= 32'hC0C0C0C1;
    10'd337 : X0 <= 32'hC09C7F27;
    10'd338 : X0 <= 32'hC0784B2F;
    10'd339 : X0 <= 32'hC05424D0;
    10'd340 : X0 <= 32'hC0300C03;
    10'd341 : X0 <= 32'hC00C00C0;
    10'd342 : X0 <= 32'hBFE80300;
    10'd343 : X0 <= 32'hBFC412BA;
    10'd344 : X0 <= 32'hBFA02FE8;
    10'd345 : X0 <= 32'hBF7C5A82;
    10'd346 : X0 <= 32'hBF589280;
    10'd347 : X0 <= 32'hBF34D7DB;
    10'd348 : X0 <= 32'hBF112A8B;
    10'd349 : X0 <= 32'hBEED8A89;
    10'd350 : X0 <= 32'hBEC9F7CD;
    10'd351 : X0 <= 32'hBEA67251;
    10'd352 : X0 <= 32'hBE82FA0C;
    10'd353 : X0 <= 32'hBE5F8EF7;
    10'd354 : X0 <= 32'hBE3C310C;
    10'd355 : X0 <= 32'hBE18E041;
    10'd356 : X0 <= 32'hBDF59C91;
    10'd357 : X0 <= 32'hBDD265F5;
    10'd358 : X0 <= 32'hBDAF3C63;
    10'd359 : X0 <= 32'hBD8C1FD7;
    10'd360 : X0 <= 32'hBD691047;
    10'd361 : X0 <= 32'hBD460DAE;
    10'd362 : X0 <= 32'hBD231803;
    10'd363 : X0 <= 32'hBD002F40;
    10'd364 : X0 <= 32'hBCDD535E;
    10'd365 : X0 <= 32'hBCBA8455;
    10'd366 : X0 <= 32'hBC97C21E;
    10'd367 : X0 <= 32'hBC750CB3;
    10'd368 : X0 <= 32'hBC52640C;
    10'd369 : X0 <= 32'hBC2FC822;
    10'd370 : X0 <= 32'hBC0D38EE;
    10'd371 : X0 <= 32'hBBEAB669;
    10'd372 : X0 <= 32'hBBC8408D;
    10'd373 : X0 <= 32'hBBA5D752;
    10'd374 : X0 <= 32'hBB837AB1;
    10'd375 : X0 <= 32'hBB612AA3;
    10'd376 : X0 <= 32'hBB3EE722;
    10'd377 : X0 <= 32'hBB1CB026;
    10'd378 : X0 <= 32'hBAFA85A9;
    10'd379 : X0 <= 32'hBAD867A4;
    10'd380 : X0 <= 32'hBAB65610;
    10'd381 : X0 <= 32'hBA9450E6;
    10'd382 : X0 <= 32'hBA725820;
    10'd383 : X0 <= 32'hBA506BB6;
    10'd384 : X0 <= 32'hBA2E8BA3;
    10'd385 : X0 <= 32'hBA0CB7DF;
    10'd386 : X0 <= 32'hB9EAF063;
    10'd387 : X0 <= 32'hB9C93529;
    10'd388 : X0 <= 32'hB9A7862A;
    10'd389 : X0 <= 32'hB985E360;
    10'd390 : X0 <= 32'hB9644CC4;
    10'd391 : X0 <= 32'hB942C24F;
    10'd392 : X0 <= 32'hB92143FA;
    10'd393 : X0 <= 32'hB8FFD1C0;
    10'd394 : X0 <= 32'hB8DE6B99;
    10'd395 : X0 <= 32'hB8BD1180;
    10'd396 : X0 <= 32'hB89BC36D;
    10'd397 : X0 <= 32'hB87A815A;
    10'd398 : X0 <= 32'hB8594B40;
    10'd399 : X0 <= 32'hB838211A;
    10'd400 : X0 <= 32'hB81702E0;
    10'd401 : X0 <= 32'hB7F5F08D;
    10'd402 : X0 <= 32'hB7D4EA19;
    10'd403 : X0 <= 32'hB7B3EF7F;
    10'd404 : X0 <= 32'hB79300B8;
    10'd405 : X0 <= 32'hB7721DBD;
    10'd406 : X0 <= 32'hB7514689;
    10'd407 : X0 <= 32'hB7307B15;
    10'd408 : X0 <= 32'hB70FBB5A;
    10'd409 : X0 <= 32'hB6EF0753;
    10'd410 : X0 <= 32'hB6CE5EF9;
    10'd411 : X0 <= 32'hB6ADC246;
    10'd412 : X0 <= 32'hB68D3134;
    10'd413 : X0 <= 32'hB66CABBC;
    10'd414 : X0 <= 32'hB64C31D9;
    10'd415 : X0 <= 32'hB62BC383;
    10'd416 : X0 <= 32'hB60B60B6;
    10'd417 : X0 <= 32'hB5EB096A;
    10'd418 : X0 <= 32'hB5CABD9A;
    10'd419 : X0 <= 32'hB5AA7D40;
    10'd420 : X0 <= 32'hB58A4855;
    10'd421 : X0 <= 32'hB56A1ED4;
    10'd422 : X0 <= 32'hB54A00B5;
    10'd423 : X0 <= 32'hB529EDF4;
    10'd424 : X0 <= 32'hB509E68B;
    10'd425 : X0 <= 32'hB4E9EA72;
    10'd426 : X0 <= 32'hB4C9F9A5;
    10'd427 : X0 <= 32'hB4AA141D;
    10'd428 : X0 <= 32'hB48A39D4;
    10'd429 : X0 <= 32'hB46A6AC5;
    10'd430 : X0 <= 32'hB44AA6E9;
    10'd431 : X0 <= 32'hB42AEE3B;
    10'd432 : X0 <= 32'hB40B40B4;
    10'd433 : X0 <= 32'hB3EB9E4F;
    10'd434 : X0 <= 32'hB3CC0706;
    10'd435 : X0 <= 32'hB3AC7AD3;
    10'd436 : X0 <= 32'hB38CF9B0;
    10'd437 : X0 <= 32'hB36D8398;
    10'd438 : X0 <= 32'hB34E1884;
    10'd439 : X0 <= 32'hB32EB86F;
    10'd440 : X0 <= 32'hB30F6353;
    10'd441 : X0 <= 32'hB2F0192A;
    10'd442 : X0 <= 32'hB2D0D9EF;
    10'd443 : X0 <= 32'hB2B1A59B;
    10'd444 : X0 <= 32'hB2927C2A;
    10'd445 : X0 <= 32'hB2735D95;
    10'd446 : X0 <= 32'hB25449D7;
    10'd447 : X0 <= 32'hB23540EA;
    10'd448 : X0 <= 32'hB21642C8;
    10'd449 : X0 <= 32'hB1F74F6D;
    10'd450 : X0 <= 32'hB1D866D1;
    10'd451 : X0 <= 32'hB1B988F0;
    10'd452 : X0 <= 32'hB19AB5C4;
    10'd453 : X0 <= 32'hB17BED48;
    10'd454 : X0 <= 32'hB15D2F75;
    10'd455 : X0 <= 32'hB13E7C47;
    10'd456 : X0 <= 32'hB11FD3B8;
    10'd457 : X0 <= 32'hB10135C2;
    10'd458 : X0 <= 32'hB0E2A260;
    10'd459 : X0 <= 32'hB0C4198C;
    10'd460 : X0 <= 32'hB0A59B42;
    10'd461 : X0 <= 32'hB087277A;
    10'd462 : X0 <= 32'hB068BE31;
    10'd463 : X0 <= 32'hB04A5F60;
    10'd464 : X0 <= 32'hB02C0B03;
    10'd465 : X0 <= 32'hB00DC113;
    10'd466 : X0 <= 32'hAFEF818C;
    10'd467 : X0 <= 32'hAFD14C68;
    10'd468 : X0 <= 32'hAFB321A1;
    10'd469 : X0 <= 32'hAF950133;
    10'd470 : X0 <= 32'hAF76EB18;
    10'd471 : X0 <= 32'hAF58DF4B;
    10'd472 : X0 <= 32'hAF3ADDC7;
    10'd473 : X0 <= 32'hAF1CE685;
    10'd474 : X0 <= 32'hAEFEF982;
    10'd475 : X0 <= 32'hAEE116B7;
    10'd476 : X0 <= 32'hAEC33E1F;
    10'd477 : X0 <= 32'hAEA56FB6;
    10'd478 : X0 <= 32'hAE87AB76;
    10'd479 : X0 <= 32'hAE69F15A;
    10'd480 : X0 <= 32'hAE4C415D;
    10'd481 : X0 <= 32'hAE2E9B79;
    10'd482 : X0 <= 32'hAE10FFA9;
    10'd483 : X0 <= 32'hADF36DE9;
    10'd484 : X0 <= 32'hADD5E632;
    10'd485 : X0 <= 32'hADB86881;
    10'd486 : X0 <= 32'hAD9AF4D0;
    10'd487 : X0 <= 32'hAD7D8B19;
    10'd488 : X0 <= 32'hAD602B58;
    10'd489 : X0 <= 32'hAD42D588;
    10'd490 : X0 <= 32'hAD2589A3;
    10'd491 : X0 <= 32'hAD0847A5;
    10'd492 : X0 <= 32'hACEB0F89;
    10'd493 : X0 <= 32'hACCDE149;
    10'd494 : X0 <= 32'hACB0BCE1;
    10'd495 : X0 <= 32'hAC93A24C;
    10'd496 : X0 <= 32'hAC769184;
    10'd497 : X0 <= 32'hAC598A85;
    10'd498 : X0 <= 32'hAC3C8D4A;
    10'd499 : X0 <= 32'hAC1F99CD;
    10'd500 : X0 <= 32'hAC02B00B;
    10'd501 : X0 <= 32'hABE5CFFD;
    10'd502 : X0 <= 32'hABC8F9A0;
    10'd503 : X0 <= 32'hABAC2CEE;
    10'd504 : X0 <= 32'hAB8F69E3;
    10'd505 : X0 <= 32'hAB72B079;
    10'd506 : X0 <= 32'hAB5600AB;
    10'd507 : X0 <= 32'hAB395A76;
    10'd508 : X0 <= 32'hAB1CBDD4;
    10'd509 : X0 <= 32'hAB002AC0;
    10'd510 : X0 <= 32'hAAE3A136;
    10'd511 : X0 <= 32'hAAC72130;
    10'd512 : X0 <= 32'hAAAAAAAB;
    10'd513 : X0 <= 32'hAA8E3DA0;
    10'd514 : X0 <= 32'hAA71DA0D;
    10'd515 : X0 <= 32'hAA557FEB;
    10'd516 : X0 <= 32'hAA392F36;
    10'd517 : X0 <= 32'hAA1CE7E9;
    10'd518 : X0 <= 32'hAA00AA01;
    10'd519 : X0 <= 32'hA9E47577;
    10'd520 : X0 <= 32'hA9C84A48;
    10'd521 : X0 <= 32'hA9AC286E;
    10'd522 : X0 <= 32'hA9900FE6;
    10'd523 : X0 <= 32'hA97400A9;
    10'd524 : X0 <= 32'hA957FAB5;
    10'd525 : X0 <= 32'hA93BFE04;
    10'd526 : X0 <= 32'hA9200A92;
    10'd527 : X0 <= 32'hA904205A;
    10'd528 : X0 <= 32'hA8E83F57;
    10'd529 : X0 <= 32'hA8CC6785;
    10'd530 : X0 <= 32'hA8B098E0;
    10'd531 : X0 <= 32'hA894D363;
    10'd532 : X0 <= 32'hA8791709;
    10'd533 : X0 <= 32'hA85D63CD;
    10'd534 : X0 <= 32'hA841B9AD;
    10'd535 : X0 <= 32'hA82618A2;
    10'd536 : X0 <= 32'hA80A80A8;
    10'd537 : X0 <= 32'hA7EEF1BB;
    10'd538 : X0 <= 32'hA7D36BD7;
    10'd539 : X0 <= 32'hA7B7EEF7;
    10'd540 : X0 <= 32'hA79C7B17;
    10'd541 : X0 <= 32'hA7811032;
    10'd542 : X0 <= 32'hA765AE43;
    10'd543 : X0 <= 32'hA74A5547;
    10'd544 : X0 <= 32'hA72F0539;
    10'd545 : X0 <= 32'hA713BE15;
    10'd546 : X0 <= 32'hA6F87FD6;
    10'd547 : X0 <= 32'hA6DD4A78;
    10'd548 : X0 <= 32'hA6C21DF7;
    10'd549 : X0 <= 32'hA6A6FA4E;
    10'd550 : X0 <= 32'hA68BDF79;
    10'd551 : X0 <= 32'hA670CD73;
    10'd552 : X0 <= 32'hA655C439;
    10'd553 : X0 <= 32'hA63AC3C6;
    10'd554 : X0 <= 32'hA61FCC16;
    10'd555 : X0 <= 32'hA604DD24;
    10'd556 : X0 <= 32'hA5E9F6ED;
    10'd557 : X0 <= 32'hA5CF196C;
    10'd558 : X0 <= 32'hA5B4449D;
    10'd559 : X0 <= 32'hA599787B;
    10'd560 : X0 <= 32'hA57EB503;
    10'd561 : X0 <= 32'hA563FA2F;
    10'd562 : X0 <= 32'hA54947FD;
    10'd563 : X0 <= 32'hA52E9E68;
    10'd564 : X0 <= 32'hA513FD6C;
    10'd565 : X0 <= 32'hA4F96504;
    10'd566 : X0 <= 32'hA4DED52C;
    10'd567 : X0 <= 32'hA4C44DE1;
    10'd568 : X0 <= 32'hA4A9CF1E;
    10'd569 : X0 <= 32'hA48F58DE;
    10'd570 : X0 <= 32'hA474EB1F;
    10'd571 : X0 <= 32'hA45A85DC;
    10'd572 : X0 <= 32'hA4402910;
    10'd573 : X0 <= 32'hA425D4B8;
    10'd574 : X0 <= 32'hA40B88D0;
    10'd575 : X0 <= 32'hA3F14553;
    10'd576 : X0 <= 32'hA3D70A3D;
    10'd577 : X0 <= 32'hA3BCD78C;
    10'd578 : X0 <= 32'hA3A2AD39;
    10'd579 : X0 <= 32'hA3888B42;
    10'd580 : X0 <= 32'hA36E71A3;
    10'd581 : X0 <= 32'hA3546057;
    10'd582 : X0 <= 32'hA33A575A;
    10'd583 : X0 <= 32'hA32056A9;
    10'd584 : X0 <= 32'hA3065E40;
    10'd585 : X0 <= 32'hA2EC6E1A;
    10'd586 : X0 <= 32'hA2D28634;
    10'd587 : X0 <= 32'hA2B8A689;
    10'd588 : X0 <= 32'hA29ECF16;
    10'd589 : X0 <= 32'hA284FFD7;
    10'd590 : X0 <= 32'hA26B38C8;
    10'd591 : X0 <= 32'hA25179E6;
    10'd592 : X0 <= 32'hA237C32B;
    10'd593 : X0 <= 32'hA21E1495;
    10'd594 : X0 <= 32'hA2046E1F;
    10'd595 : X0 <= 32'hA1EACFC6;
    10'd596 : X0 <= 32'hA1D13985;
    10'd597 : X0 <= 32'hA1B7AB5A;
    10'd598 : X0 <= 32'hA19E253F;
    10'd599 : X0 <= 32'hA184A732;
    10'd600 : X0 <= 32'hA16B312F;
    10'd601 : X0 <= 32'hA151C331;
    10'd602 : X0 <= 32'hA1385D35;
    10'd603 : X0 <= 32'hA11EFF37;
    10'd604 : X0 <= 32'hA105A933;
    10'd605 : X0 <= 32'hA0EC5B26;
    10'd606 : X0 <= 32'hA0D3150C;
    10'd607 : X0 <= 32'hA0B9D6E0;
    10'd608 : X0 <= 32'hA0A0A0A1;
    10'd609 : X0 <= 32'hA0877248;
    10'd610 : X0 <= 32'hA06E4BD4;
    10'd611 : X0 <= 32'hA0552D40;
    10'd612 : X0 <= 32'hA03C1688;
    10'd613 : X0 <= 32'hA02307AA;
    10'd614 : X0 <= 32'hA00A00A0;
    10'd615 : X0 <= 32'h9FF10168;
    10'd616 : X0 <= 32'h9FD809FE;
    10'd617 : X0 <= 32'h9FBF1A5D;
    10'd618 : X0 <= 32'h9FA63284;
    10'd619 : X0 <= 32'h9F8D526D;
    10'd620 : X0 <= 32'h9F747A15;
    10'd621 : X0 <= 32'h9F5BA979;
    10'd622 : X0 <= 32'h9F42E095;
    10'd623 : X0 <= 32'h9F2A1F66;
    10'd624 : X0 <= 32'h9F1165E7;
    10'd625 : X0 <= 32'h9EF8B416;
    10'd626 : X0 <= 32'h9EE009EE;
    10'd627 : X0 <= 32'h9EC7676C;
    10'd628 : X0 <= 32'h9EAECC8D;
    10'd629 : X0 <= 32'h9E96394D;
    10'd630 : X0 <= 32'h9E7DADA9;
    10'd631 : X0 <= 32'h9E65299C;
    10'd632 : X0 <= 32'h9E4CAD24;
    10'd633 : X0 <= 32'h9E34383D;
    10'd634 : X0 <= 32'h9E1BCAE3;
    10'd635 : X0 <= 32'h9E036513;
    10'd636 : X0 <= 32'h9DEB06C9;
    10'd637 : X0 <= 32'h9DD2B002;
    10'd638 : X0 <= 32'h9DBA60BB;
    10'd639 : X0 <= 32'h9DA218F0;
    10'd640 : X0 <= 32'h9D89D89E;
    10'd641 : X0 <= 32'h9D719FC0;
    10'd642 : X0 <= 32'h9D596E54;
    10'd643 : X0 <= 32'h9D414457;
    10'd644 : X0 <= 32'h9D2921C4;
    10'd645 : X0 <= 32'h9D110698;
    10'd646 : X0 <= 32'h9CF8F2D1;
    10'd647 : X0 <= 32'h9CE0E66A;
    10'd648 : X0 <= 32'h9CC8E161;
    10'd649 : X0 <= 32'h9CB0E3B1;
    10'd650 : X0 <= 32'h9C98ED58;
    10'd651 : X0 <= 32'h9C80FE52;
    10'd652 : X0 <= 32'h9C69169B;
    10'd653 : X0 <= 32'h9C513631;
    10'd654 : X0 <= 32'h9C395D10;
    10'd655 : X0 <= 32'h9C218B35;
    10'd656 : X0 <= 32'h9C09C09C;
    10'd657 : X0 <= 32'h9BF1FD42;
    10'd658 : X0 <= 32'h9BDA4124;
    10'd659 : X0 <= 32'h9BC28C3F;
    10'd660 : X0 <= 32'h9BAADE8E;
    10'd661 : X0 <= 32'h9B933810;
    10'd662 : X0 <= 32'h9B7B98C0;
    10'd663 : X0 <= 32'h9B64009B;
    10'd664 : X0 <= 32'h9B4C6F9F;
    10'd665 : X0 <= 32'h9B34E5C7;
    10'd666 : X0 <= 32'h9B1D6311;
    10'd667 : X0 <= 32'h9B05E77A;
    10'd668 : X0 <= 32'h9AEE72FD;
    10'd669 : X0 <= 32'h9AD70598;
    10'd670 : X0 <= 32'h9ABF9F48;
    10'd671 : X0 <= 32'h9AA8400A;
    10'd672 : X0 <= 32'h9A90E7D9;
    10'd673 : X0 <= 32'h9A7996B4;
    10'd674 : X0 <= 32'h9A624C97;
    10'd675 : X0 <= 32'h9A4B097E;
    10'd676 : X0 <= 32'h9A33CD67;
    10'd677 : X0 <= 32'h9A1C984E;
    10'd678 : X0 <= 32'h9A056A31;
    10'd679 : X0 <= 32'h99EE430B;
    10'd680 : X0 <= 32'h99D722DB;
    10'd681 : X0 <= 32'h99C0099C;
    10'd682 : X0 <= 32'h99A8F74C;
    10'd683 : X0 <= 32'h9991EBE7;
    10'd684 : X0 <= 32'h997AE76B;
    10'd685 : X0 <= 32'h9963E9D5;
    10'd686 : X0 <= 32'h994CF320;
    10'd687 : X0 <= 32'h9936034B;
    10'd688 : X0 <= 32'h991F1A51;
    10'd689 : X0 <= 32'h99083831;
    10'd690 : X0 <= 32'h98F15CE7;
    10'd691 : X0 <= 32'h98DA886F;
    10'd692 : X0 <= 32'h98C3BAC7;
    10'd693 : X0 <= 32'h98ACF3EC;
    10'd694 : X0 <= 32'h989633DB;
    10'd695 : X0 <= 32'h987F7A90;
    10'd696 : X0 <= 32'h9868C80A;
    10'd697 : X0 <= 32'h98521C43;
    10'd698 : X0 <= 32'h983B773B;
    10'd699 : X0 <= 32'h9824D8ED;
    10'd700 : X0 <= 32'h980E4156;
    10'd701 : X0 <= 32'h97F7B074;
    10'd702 : X0 <= 32'h97E12644;
    10'd703 : X0 <= 32'h97CAA2C3;
    10'd704 : X0 <= 32'h97B425ED;
    10'd705 : X0 <= 32'h979DAFC0;
    10'd706 : X0 <= 32'h97874039;
    10'd707 : X0 <= 32'h9770D754;
    10'd708 : X0 <= 32'h975A7510;
    10'd709 : X0 <= 32'h97441968;
    10'd710 : X0 <= 32'h972DC45B;
    10'd711 : X0 <= 32'h971775E5;
    10'd712 : X0 <= 32'h97012E02;
    10'd713 : X0 <= 32'h96EAECB1;
    10'd714 : X0 <= 32'h96D4B1EF;
    10'd715 : X0 <= 32'h96BE7DB8;
    10'd716 : X0 <= 32'h96A85009;
    10'd717 : X0 <= 32'h969228E1;
    10'd718 : X0 <= 32'h967C083B;
    10'd719 : X0 <= 32'h9665EE15;
    10'd720 : X0 <= 32'h964FDA6C;
    10'd721 : X0 <= 32'h9639CD3D;
    10'd722 : X0 <= 32'h9623C686;
    10'd723 : X0 <= 32'h960DC644;
    10'd724 : X0 <= 32'h95F7CC73;
    10'd725 : X0 <= 32'h95E1D911;
    10'd726 : X0 <= 32'h95CBEC1B;
    10'd727 : X0 <= 32'h95B6058E;
    10'd728 : X0 <= 32'h95A02568;
    10'd729 : X0 <= 32'h958A4BA5;
    10'd730 : X0 <= 32'h95747844;
    10'd731 : X0 <= 32'h955EAB40;
    10'd732 : X0 <= 32'h9548E498;
    10'd733 : X0 <= 32'h95332448;
    10'd734 : X0 <= 32'h951D6A4D;
    10'd735 : X0 <= 32'h9507B6A6;
    10'd736 : X0 <= 32'h94F2094F;
    10'd737 : X0 <= 32'h94DC6245;
    10'd738 : X0 <= 32'h94C6C187;
    10'd739 : X0 <= 32'h94B12710;
    10'd740 : X0 <= 32'h949B92DE;
    10'd741 : X0 <= 32'h948604EE;
    10'd742 : X0 <= 32'h94707D3F;
    10'd743 : X0 <= 32'h945AFBCC;
    10'd744 : X0 <= 32'h94458094;
    10'd745 : X0 <= 32'h94300B94;
    10'd746 : X0 <= 32'h941A9CC8;
    10'd747 : X0 <= 32'h9405342F;
    10'd748 : X0 <= 32'h93EFD1C5;
    10'd749 : X0 <= 32'h93DA7588;
    10'd750 : X0 <= 32'h93C51F75;
    10'd751 : X0 <= 32'h93AFCF8A;
    10'd752 : X0 <= 32'h939A85C4;
    10'd753 : X0 <= 32'h93854220;
    10'd754 : X0 <= 32'h9370049C;
    10'd755 : X0 <= 32'h935ACD34;
    10'd756 : X0 <= 32'h93459BE7;
    10'd757 : X0 <= 32'h933070B1;
    10'd758 : X0 <= 32'h931B4B91;
    10'd759 : X0 <= 32'h93062C82;
    10'd760 : X0 <= 32'h92F11384;
    10'd761 : X0 <= 32'h92DC0093;
    10'd762 : X0 <= 32'h92C6F3AC;
    10'd763 : X0 <= 32'h92B1ECCE;
    10'd764 : X0 <= 32'h929CEBF5;
    10'd765 : X0 <= 32'h9287F11E;
    10'd766 : X0 <= 32'h9272FC48;
    10'd767 : X0 <= 32'h925E0D70;
    10'd768 : X0 <= 32'h92492492;
    10'd769 : X0 <= 32'h923441AD;
    10'd770 : X0 <= 32'h921F64BF;
    10'd771 : X0 <= 32'h920A8DC3;
    10'd772 : X0 <= 32'h91F5BCB9;
    10'd773 : X0 <= 32'h91E0F19D;
    10'd774 : X0 <= 32'h91CC2C6C;
    10'd775 : X0 <= 32'h91B76D25;
    10'd776 : X0 <= 32'h91A2B3C5;
    10'd777 : X0 <= 32'h918E0049;
    10'd778 : X0 <= 32'h917952AE;
    10'd779 : X0 <= 32'h9164AAF3;
    10'd780 : X0 <= 32'h91500915;
    10'd781 : X0 <= 32'h913B6D11;
    10'd782 : X0 <= 32'h9126D6E5;
    10'd783 : X0 <= 32'h9112468D;
    10'd784 : X0 <= 32'h90FDBC09;
    10'd785 : X0 <= 32'h90E93755;
    10'd786 : X0 <= 32'h90D4B86F;
    10'd787 : X0 <= 32'h90C03F54;
    10'd788 : X0 <= 32'h90ABCC02;
    10'd789 : X0 <= 32'h90975E77;
    10'd790 : X0 <= 32'h9082F6B0;
    10'd791 : X0 <= 32'h906E94AA;
    10'd792 : X0 <= 32'h905A3863;
    10'd793 : X0 <= 32'h9045E1D9;
    10'd794 : X0 <= 32'h9031910A;
    10'd795 : X0 <= 32'h901D45F2;
    10'd796 : X0 <= 32'h90090090;
    10'd797 : X0 <= 32'h8FF4C0E1;
    10'd798 : X0 <= 32'h8FE086E2;
    10'd799 : X0 <= 32'h8FCC5292;
    10'd800 : X0 <= 32'h8FB823EE;
    10'd801 : X0 <= 32'h8FA3FAF3;
    10'd802 : X0 <= 32'h8F8FD7A0;
    10'd803 : X0 <= 32'h8F7BB9F1;
    10'd804 : X0 <= 32'h8F67A1E4;
    10'd805 : X0 <= 32'h8F538F77;
    10'd806 : X0 <= 32'h8F3F82A8;
    10'd807 : X0 <= 32'h8F2B7B75;
    10'd808 : X0 <= 32'h8F1779DA;
    10'd809 : X0 <= 32'h8F037DD6;
    10'd810 : X0 <= 32'h8EEF8766;
    10'd811 : X0 <= 32'h8EDB9688;
    10'd812 : X0 <= 32'h8EC7AB39;
    10'd813 : X0 <= 32'h8EB3C578;
    10'd814 : X0 <= 32'h8E9FE542;
    10'd815 : X0 <= 32'h8E8C0A94;
    10'd816 : X0 <= 32'h8E78356D;
    10'd817 : X0 <= 32'h8E6465CA;
    10'd818 : X0 <= 32'h8E509BA8;
    10'd819 : X0 <= 32'h8E3CD706;
    10'd820 : X0 <= 32'h8E2917E1;
    10'd821 : X0 <= 32'h8E155E37;
    10'd822 : X0 <= 32'h8E01AA05;
    10'd823 : X0 <= 32'h8DEDFB4A;
    10'd824 : X0 <= 32'h8DDA5202;
    10'd825 : X0 <= 32'h8DC6AE2D;
    10'd826 : X0 <= 32'h8DB30FC6;
    10'd827 : X0 <= 32'h8D9F76CE;
    10'd828 : X0 <= 32'h8D8BE340;
    10'd829 : X0 <= 32'h8D78551A;
    10'd830 : X0 <= 32'h8D64CC5C;
    10'd831 : X0 <= 32'h8D514901;
    10'd832 : X0 <= 32'h8D3DCB09;
    10'd833 : X0 <= 32'h8D2A5270;
    10'd834 : X0 <= 32'h8D16DF35;
    10'd835 : X0 <= 32'h8D037156;
    10'd836 : X0 <= 32'h8CF008CF;
    10'd837 : X0 <= 32'h8CDCA59F;
    10'd838 : X0 <= 32'h8CC947C5;
    10'd839 : X0 <= 32'h8CB5EF3C;
    10'd840 : X0 <= 32'h8CA29C04;
    10'd841 : X0 <= 32'h8C8F4E1B;
    10'd842 : X0 <= 32'h8C7C057D;
    10'd843 : X0 <= 32'h8C68C229;
    10'd844 : X0 <= 32'h8C55841D;
    10'd845 : X0 <= 32'h8C424B56;
    10'd846 : X0 <= 32'h8C2F17D2;
    10'd847 : X0 <= 32'h8C1BE990;
    10'd848 : X0 <= 32'h8C08C08C;
    10'd849 : X0 <= 32'h8BF59CC5;
    10'd850 : X0 <= 32'h8BE27E39;
    10'd851 : X0 <= 32'h8BCF64E6;
    10'd852 : X0 <= 32'h8BBC50C9;
    10'd853 : X0 <= 32'h8BA941E0;
    10'd854 : X0 <= 32'h8B963829;
    10'd855 : X0 <= 32'h8B8333A3;
    10'd856 : X0 <= 32'h8B70344A;
    10'd857 : X0 <= 32'h8B5D3A1D;
    10'd858 : X0 <= 32'h8B4A451A;
    10'd859 : X0 <= 32'h8B37553E;
    10'd860 : X0 <= 32'h8B246A88;
    10'd861 : X0 <= 32'h8B1184F5;
    10'd862 : X0 <= 32'h8AFEA483;
    10'd863 : X0 <= 32'h8AEBC931;
    10'd864 : X0 <= 32'h8AD8F2FC;
    10'd865 : X0 <= 32'h8AC621E1;
    10'd866 : X0 <= 32'h8AB355E0;
    10'd867 : X0 <= 32'h8AA08EF6;
    10'd868 : X0 <= 32'h8A8DCD20;
    10'd869 : X0 <= 32'h8A7B105D;
    10'd870 : X0 <= 32'h8A6858AB;
    10'd871 : X0 <= 32'h8A55A607;
    10'd872 : X0 <= 32'h8A42F870;
    10'd873 : X0 <= 32'h8A304FE4;
    10'd874 : X0 <= 32'h8A1DAC60;
    10'd875 : X0 <= 32'h8A0B0DE3;
    10'd876 : X0 <= 32'h89F8746A;
    10'd877 : X0 <= 32'h89E5DFF3;
    10'd878 : X0 <= 32'h89D3507D;
    10'd879 : X0 <= 32'h89C0C605;
    10'd880 : X0 <= 32'h89AE408A;
    10'd881 : X0 <= 32'h899BC009;
    10'd882 : X0 <= 32'h89894480;
    10'd883 : X0 <= 32'h8976CDED;
    10'd884 : X0 <= 32'h89645C4F;
    10'd885 : X0 <= 32'h8951EFA4;
    10'd886 : X0 <= 32'h893F87E8;
    10'd887 : X0 <= 32'h892D251B;
    10'd888 : X0 <= 32'h891AC73B;
    10'd889 : X0 <= 32'h89086E45;
    10'd890 : X0 <= 32'h88F61A37;
    10'd891 : X0 <= 32'h88E3CB10;
    10'd892 : X0 <= 32'h88D180CD;
    10'd893 : X0 <= 32'h88BF3B6D;
    10'd894 : X0 <= 32'h88ACFAEE;
    10'd895 : X0 <= 32'h889ABF4D;
    10'd896 : X0 <= 32'h88888889;
    10'd897 : X0 <= 32'h8876569F;
    10'd898 : X0 <= 32'h8864298F;
    10'd899 : X0 <= 32'h88520155;
    10'd900 : X0 <= 32'h883FDDF0;
    10'd901 : X0 <= 32'h882DBF5E;
    10'd902 : X0 <= 32'h881BA59E;
    10'd903 : X0 <= 32'h880990AC;
    10'd904 : X0 <= 32'h87F78088;
    10'd905 : X0 <= 32'h87E5752F;
    10'd906 : X0 <= 32'h87D36EA0;
    10'd907 : X0 <= 32'h87C16CD8;
    10'd908 : X0 <= 32'h87AF6FD6;
    10'd909 : X0 <= 32'h879D7797;
    10'd910 : X0 <= 32'h878B841A;
    10'd911 : X0 <= 32'h8779955E;
    10'd912 : X0 <= 32'h8767AB5F;
    10'd913 : X0 <= 32'h8755C61D;
    10'd914 : X0 <= 32'h8743E595;
    10'd915 : X0 <= 32'h873209C5;
    10'd916 : X0 <= 32'h872032AC;
    10'd917 : X0 <= 32'h870E6048;
    10'd918 : X0 <= 32'h86FC9296;
    10'd919 : X0 <= 32'h86EAC996;
    10'd920 : X0 <= 32'h86D90544;
    10'd921 : X0 <= 32'h86C745A0;
    10'd922 : X0 <= 32'h86B58AA8;
    10'd923 : X0 <= 32'h86A3D459;
    10'd924 : X0 <= 32'h869222B2;
    10'd925 : X0 <= 32'h868075B0;
    10'd926 : X0 <= 32'h866ECD53;
    10'd927 : X0 <= 32'h865D2998;
    10'd928 : X0 <= 32'h864B8A7E;
    10'd929 : X0 <= 32'h8639F002;
    10'd930 : X0 <= 32'h86285A23;
    10'd931 : X0 <= 32'h8616C8DF;
    10'd932 : X0 <= 32'h86053C34;
    10'd933 : X0 <= 32'h85F3B421;
    10'd934 : X0 <= 32'h85E230A3;
    10'd935 : X0 <= 32'h85D0B1B9;
    10'd936 : X0 <= 32'h85BF3761;
    10'd937 : X0 <= 32'h85ADC199;
    10'd938 : X0 <= 32'h859C5060;
    10'd939 : X0 <= 32'h858AE3B3;
    10'd940 : X0 <= 32'h85797B91;
    10'd941 : X0 <= 32'h856817F9;
    10'd942 : X0 <= 32'h8556B8E7;
    10'd943 : X0 <= 32'h85455E5B;
    10'd944 : X0 <= 32'h85340853;
    10'd945 : X0 <= 32'h8522B6CD;
    10'd946 : X0 <= 32'h851169C7;
    10'd947 : X0 <= 32'h85002140;
    10'd948 : X0 <= 32'h84EEDD35;
    10'd949 : X0 <= 32'h84DD9DA6;
    10'd950 : X0 <= 32'h84CC6290;
    10'd951 : X0 <= 32'h84BB2BF1;
    10'd952 : X0 <= 32'h84A9F9C8;
    10'd953 : X0 <= 32'h8498CC13;
    10'd954 : X0 <= 32'h8487A2D1;
    10'd955 : X0 <= 32'h84767DFF;
    10'd956 : X0 <= 32'h84655D9C;
    10'd957 : X0 <= 32'h845441A6;
    10'd958 : X0 <= 32'h84432A1B;
    10'd959 : X0 <= 32'h843216FB;
    10'd960 : X0 <= 32'h84210842;
    10'd961 : X0 <= 32'h840FFDF0;
    10'd962 : X0 <= 32'h83FEF802;
    10'd963 : X0 <= 32'h83EDF677;
    10'd964 : X0 <= 32'h83DCF94E;
    10'd965 : X0 <= 32'h83CC0084;
    10'd966 : X0 <= 32'h83BB0C18;
    10'd967 : X0 <= 32'h83AA1C08;
    10'd968 : X0 <= 32'h83993052;
    10'd969 : X0 <= 32'h838848F6;
    10'd970 : X0 <= 32'h837765F0;
    10'd971 : X0 <= 32'h83668740;
    10'd972 : X0 <= 32'h8355ACE4;
    10'd973 : X0 <= 32'h8344D6DA;
    10'd974 : X0 <= 32'h83340520;
    10'd975 : X0 <= 32'h832337B5;
    10'd976 : X0 <= 32'h83126E98;
    10'd977 : X0 <= 32'h8301A9C5;
    10'd978 : X0 <= 32'h82F0E93D;
    10'd979 : X0 <= 32'h82E02CFD;
    10'd980 : X0 <= 32'h82CF7504;
    10'd981 : X0 <= 32'h82BEC14F;
    10'd982 : X0 <= 32'h82AE11DE;
    10'd983 : X0 <= 32'h829D66AE;
    10'd984 : X0 <= 32'h828CBFBF;
    10'd985 : X0 <= 32'h827C1D0E;
    10'd986 : X0 <= 32'h826B7E99;
    10'd987 : X0 <= 32'h825AE460;
    10'd988 : X0 <= 32'h824A4E61;
    10'd989 : X0 <= 32'h8239BC99;
    10'd990 : X0 <= 32'h82292F08;
    10'd991 : X0 <= 32'h8218A5AB;
    10'd992 : X0 <= 32'h82082082;
    10'd993 : X0 <= 32'h81F79F8A;
    10'd994 : X0 <= 32'h81E722C2;
    10'd995 : X0 <= 32'h81D6AA29;
    10'd996 : X0 <= 32'h81C635BC;
    10'd997 : X0 <= 32'h81B5C57A;
    10'd998 : X0 <= 32'h81A55963;
    10'd999 : X0 <= 32'h8194F173;
    10'd1000 : X0 <= 32'h81848DA9;
    10'd1001 : X0 <= 32'h81742E04;
    10'd1002 : X0 <= 32'h8163D283;
    10'd1003 : X0 <= 32'h81537B23;
    10'd1004 : X0 <= 32'h814327E4;
    10'd1005 : X0 <= 32'h8132D8C3;
    10'd1006 : X0 <= 32'h81228DBF;
    10'd1007 : X0 <= 32'h811246D7;
    10'd1008 : X0 <= 32'h81020408;
    10'd1009 : X0 <= 32'h80F1C552;
    10'd1010 : X0 <= 32'h80E18AB3;
    10'd1011 : X0 <= 32'h80D15429;
    10'd1012 : X0 <= 32'h80C121B3;
    10'd1013 : X0 <= 32'h80B0F34F;
    10'd1014 : X0 <= 32'h80A0C8FB;
    10'd1015 : X0 <= 32'h8090A2B7;
    10'd1016 : X0 <= 32'h80808081;
    10'd1017 : X0 <= 32'h80706256;
    10'd1018 : X0 <= 32'h80604836;
    10'd1019 : X0 <= 32'h8050321F;
    10'd1020 : X0 <= 32'h80402010;
    10'd1021 : X0 <= 32'h80301207;
    10'd1022 : X0 <= 32'h80200802;
    10'd1023 : X0 <= 32'h80100200;
    default : X0 <= 32'hFFFFFFFF;
  endcase
end


endmodule
